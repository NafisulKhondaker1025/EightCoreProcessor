`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/23/2021 03:13:04 PM
// Design Name: 
// Module Name: DataMemory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module DataMemory(Address, WriteData, Clk, MemWrite, MemRead, ReadData); 

    input [31:0] Address; 	                                 // Input Address 
    input [31:0] WriteData;                                  // Data that needs to be written into the address 
    input Clk;
    input MemWrite; 		                                 // Control signal for memory write 
    input MemRead; 			                                 // Control signal for memory read 
    
    output reg[31:0] ReadData;                               // Contents of memory location at Address

    reg [31:0] memory [0:8191];
    
    initial begin
    //$readmemh("data_memory.mem",memory);
    memory[0] = 32'h40;
memory[1] = 32'h40;
memory[2] = 32'h4;
memory[3] = 32'h4;
memory[4] = 32'hff;
memory[5] = 32'hfe;
memory[6] = 32'hfd;
memory[7] = 32'hfc;
memory[8] = 32'hfb;
memory[9] = 32'hfa;
memory[10] = 32'hf9;
memory[11] = 32'hf8;
memory[12] = 32'hf7;
memory[13] = 32'hf6;
memory[14] = 32'hf5;
memory[15] = 32'hf4;
memory[16] = 32'hf3;
memory[17] = 32'hf2;
memory[18] = 32'hf1;
memory[19] = 32'hf0;
memory[20] = 32'hef;
memory[21] = 32'hee;
memory[22] = 32'hed;
memory[23] = 32'hec;
memory[24] = 32'heb;
memory[25] = 32'hea;
memory[26] = 32'he9;
memory[27] = 32'he8;
memory[28] = 32'he7;
memory[29] = 32'he6;
memory[30] = 32'he5;
memory[31] = 32'he4;
memory[32] = 32'he3;
memory[33] = 32'he2;
memory[34] = 32'he1;
memory[35] = 32'hfe;
memory[36] = 32'hfd;
memory[37] = 32'hfc;
memory[38] = 32'hfb;
memory[39] = 32'hfa;
memory[40] = 32'hf9;
memory[41] = 32'hf8;
memory[42] = 32'hf7;
memory[43] = 32'hf6;
memory[44] = 32'hf5;
memory[45] = 32'hf4;
memory[46] = 32'hf3;
memory[47] = 32'hf2;
memory[48] = 32'hf1;
memory[49] = 32'hf0;
memory[50] = 32'hef;
memory[51] = 32'hee;
memory[52] = 32'hed;
memory[53] = 32'hec;
memory[54] = 32'heb;
memory[55] = 32'hea;
memory[56] = 32'he9;
memory[57] = 32'he8;
memory[58] = 32'he7;
memory[59] = 32'he6;
memory[60] = 32'he5;
memory[61] = 32'he4;
memory[62] = 32'he3;
memory[63] = 32'he2;
memory[64] = 32'he1;
memory[65] = 32'hfe;
memory[66] = 32'hfd;
memory[67] = 32'hfb;
memory[68] = 32'hf0;
memory[69] = 32'hef;
memory[70] = 32'hee;
memory[71] = 32'hed;
memory[72] = 32'hec;
memory[73] = 32'heb;
memory[74] = 32'hea;
memory[75] = 32'he9;
memory[76] = 32'he8;
memory[77] = 32'he7;
memory[78] = 32'he6;
memory[79] = 32'he5;
memory[80] = 32'he4;
memory[81] = 32'he3;
memory[82] = 32'he2;
memory[83] = 32'he1;
memory[84] = 32'hfe;
memory[85] = 32'hfd;
memory[86] = 32'hfc;
memory[87] = 32'hfb;
memory[88] = 32'hfa;
memory[89] = 32'hf9;
memory[90] = 32'hf8;
memory[91] = 32'hf7;
memory[92] = 32'hf6;
memory[93] = 32'hf5;
memory[94] = 32'hf4;
memory[95] = 32'hf3;
memory[96] = 32'hf2;
memory[97] = 32'hf1;
memory[98] = 32'hf0;
memory[99] = 32'hef;
memory[100] = 32'hee;
memory[101] = 32'hed;
memory[102] = 32'hec;
memory[103] = 32'heb;
memory[104] = 32'hea;
memory[105] = 32'he9;
memory[106] = 32'he8;
memory[107] = 32'he7;
memory[108] = 32'he6;
memory[109] = 32'he5;
memory[110] = 32'he4;
memory[111] = 32'he3;
memory[112] = 32'he2;
memory[113] = 32'he1;
memory[114] = 32'hfe;
memory[115] = 32'hfd;
memory[116] = 32'hfc;
memory[117] = 32'hfb;
memory[118] = 32'hfa;
memory[119] = 32'hf9;
memory[120] = 32'hf8;
memory[121] = 32'hf7;
memory[122] = 32'hf6;
memory[123] = 32'hf5;
memory[124] = 32'hf4;
memory[125] = 32'hf3;
memory[126] = 32'hf2;
memory[127] = 32'hf1;
memory[128] = 32'hf0;
memory[129] = 32'hef;
memory[130] = 32'hed;
memory[131] = 32'hfa;
memory[132] = 32'hf2;
memory[133] = 32'he8;
memory[134] = 32'he7;
memory[135] = 32'he6;
memory[136] = 32'he5;
memory[137] = 32'he4;
memory[138] = 32'he3;
memory[139] = 32'he2;
memory[140] = 32'he1;
memory[141] = 32'hfe;
memory[142] = 32'hfd;
memory[143] = 32'hfc;
memory[144] = 32'hfb;
memory[145] = 32'hfa;
memory[146] = 32'hf9;
memory[147] = 32'hf8;
memory[148] = 32'hf7;
memory[149] = 32'hf6;
memory[150] = 32'hf5;
memory[151] = 32'hf4;
memory[152] = 32'hf3;
memory[153] = 32'hf2;
memory[154] = 32'hf1;
memory[155] = 32'hf0;
memory[156] = 32'hef;
memory[157] = 32'hee;
memory[158] = 32'hed;
memory[159] = 32'hec;
memory[160] = 32'heb;
memory[161] = 32'hea;
memory[162] = 32'he9;
memory[163] = 32'he8;
memory[164] = 32'he7;
memory[165] = 32'he6;
memory[166] = 32'he5;
memory[167] = 32'he4;
memory[168] = 32'he3;
memory[169] = 32'he2;
memory[170] = 32'he1;
memory[171] = 32'hfe;
memory[172] = 32'hfd;
memory[173] = 32'hfc;
memory[174] = 32'hfb;
memory[175] = 32'hfa;
memory[176] = 32'hf9;
memory[177] = 32'hf8;
memory[178] = 32'hf7;
memory[179] = 32'hf6;
memory[180] = 32'hf5;
memory[181] = 32'hf4;
memory[182] = 32'hf3;
memory[183] = 32'hf2;
memory[184] = 32'hf1;
memory[185] = 32'hf0;
memory[186] = 32'hef;
memory[187] = 32'hee;
memory[188] = 32'hed;
memory[189] = 32'hec;
memory[190] = 32'heb;
memory[191] = 32'hea;
memory[192] = 32'he9;
memory[193] = 32'he7;
memory[194] = 32'hec;
memory[195] = 32'hf9;
memory[196] = 32'hf3;
memory[197] = 32'hea;
memory[198] = 32'he8;
memory[199] = 32'he7;
memory[200] = 32'he6;
memory[201] = 32'he5;
memory[202] = 32'he4;
memory[203] = 32'he3;
memory[204] = 32'he2;
memory[205] = 32'he1;
memory[206] = 32'hfe;
memory[207] = 32'hfd;
memory[208] = 32'hfc;
memory[209] = 32'hfb;
memory[210] = 32'hfa;
memory[211] = 32'hf9;
memory[212] = 32'hf8;
memory[213] = 32'hf7;
memory[214] = 32'hf6;
memory[215] = 32'hf5;
memory[216] = 32'hf4;
memory[217] = 32'hf3;
memory[218] = 32'hf2;
memory[219] = 32'hf1;
memory[220] = 32'hf0;
memory[221] = 32'hef;
memory[222] = 32'hee;
memory[223] = 32'hed;
memory[224] = 32'hec;
memory[225] = 32'heb;
memory[226] = 32'hea;
memory[227] = 32'he9;
memory[228] = 32'he8;
memory[229] = 32'he7;
memory[230] = 32'he6;
memory[231] = 32'he5;
memory[232] = 32'he4;
memory[233] = 32'he3;
memory[234] = 32'he2;
memory[235] = 32'he1;
memory[236] = 32'hfe;
memory[237] = 32'hfd;
memory[238] = 32'hfc;
memory[239] = 32'hfb;
memory[240] = 32'hfa;
memory[241] = 32'hf9;
memory[242] = 32'hf8;
memory[243] = 32'hf7;
memory[244] = 32'hf6;
memory[245] = 32'hf5;
memory[246] = 32'hf4;
memory[247] = 32'hf3;
memory[248] = 32'hf2;
memory[249] = 32'hf1;
memory[250] = 32'hf0;
memory[251] = 32'hef;
memory[252] = 32'hee;
memory[253] = 32'hed;
memory[254] = 32'hec;
memory[255] = 32'heb;
memory[256] = 32'he9;
memory[257] = 32'he6;
memory[258] = 32'heb;
memory[259] = 32'hf8;
memory[260] = 32'hf4;
memory[261] = 32'heb;
memory[262] = 32'hea;
memory[263] = 32'hf0;
memory[264] = 32'hef;
memory[265] = 32'hee;
memory[266] = 32'hed;
memory[267] = 32'hec;
memory[268] = 32'heb;
memory[269] = 32'hea;
memory[270] = 32'he9;
memory[271] = 32'he8;
memory[272] = 32'he7;
memory[273] = 32'he6;
memory[274] = 32'he5;
memory[275] = 32'he4;
memory[276] = 32'he3;
memory[277] = 32'he2;
memory[278] = 32'he1;
memory[279] = 32'hfe;
memory[280] = 32'hfd;
memory[281] = 32'hfc;
memory[282] = 32'hfb;
memory[283] = 32'hfa;
memory[284] = 32'hf9;
memory[285] = 32'hf8;
memory[286] = 32'hf7;
memory[287] = 32'hf6;
memory[288] = 32'hf5;
memory[289] = 32'hf4;
memory[290] = 32'hf3;
memory[291] = 32'hf2;
memory[292] = 32'hf1;
memory[293] = 32'hf0;
memory[294] = 32'hef;
memory[295] = 32'hee;
memory[296] = 32'hed;
memory[297] = 32'hec;
memory[298] = 32'heb;
memory[299] = 32'hea;
memory[300] = 32'he9;
memory[301] = 32'he8;
memory[302] = 32'he7;
memory[303] = 32'he6;
memory[304] = 32'he5;
memory[305] = 32'he4;
memory[306] = 32'he3;
memory[307] = 32'he2;
memory[308] = 32'he1;
memory[309] = 32'hfe;
memory[310] = 32'hfd;
memory[311] = 32'hfc;
memory[312] = 32'hfb;
memory[313] = 32'hfa;
memory[314] = 32'hf9;
memory[315] = 32'hf8;
memory[316] = 32'hf7;
memory[317] = 32'hf6;
memory[318] = 32'hf5;
memory[319] = 32'hf3;
memory[320] = 32'he8;
memory[321] = 32'he5;
memory[322] = 32'hea;
memory[323] = 32'hf7;
memory[324] = 32'hf5;
memory[325] = 32'hec;
memory[326] = 32'heb;
memory[327] = 32'hf2;
memory[328] = 32'he2;
memory[329] = 32'he1;
memory[330] = 32'hfe;
memory[331] = 32'hfd;
memory[332] = 32'hfc;
memory[333] = 32'hfb;
memory[334] = 32'hfa;
memory[335] = 32'hf9;
memory[336] = 32'hf8;
memory[337] = 32'hf7;
memory[338] = 32'hf6;
memory[339] = 32'hf5;
memory[340] = 32'hf4;
memory[341] = 32'hf3;
memory[342] = 32'hf2;
memory[343] = 32'hf1;
memory[344] = 32'hf0;
memory[345] = 32'hef;
memory[346] = 32'hee;
memory[347] = 32'hed;
memory[348] = 32'hec;
memory[349] = 32'heb;
memory[350] = 32'hea;
memory[351] = 32'he9;
memory[352] = 32'he8;
memory[353] = 32'he7;
memory[354] = 32'he6;
memory[355] = 32'he5;
memory[356] = 32'he4;
memory[357] = 32'he3;
memory[358] = 32'he2;
memory[359] = 32'he1;
memory[360] = 32'hfe;
memory[361] = 32'hfd;
memory[362] = 32'hfc;
memory[363] = 32'hfb;
memory[364] = 32'hfa;
memory[365] = 32'hf9;
memory[366] = 32'hf8;
memory[367] = 32'hf7;
memory[368] = 32'hf6;
memory[369] = 32'hf5;
memory[370] = 32'hf4;
memory[371] = 32'hf3;
memory[372] = 32'hf2;
memory[373] = 32'hf1;
memory[374] = 32'hf0;
memory[375] = 32'hef;
memory[376] = 32'hee;
memory[377] = 32'hed;
memory[378] = 32'hec;
memory[379] = 32'heb;
memory[380] = 32'hea;
memory[381] = 32'he9;
memory[382] = 32'he7;
memory[383] = 32'hf2;
memory[384] = 32'he7;
memory[385] = 32'he4;
memory[386] = 32'he9;
memory[387] = 32'hf6;
memory[388] = 32'hf6;
memory[389] = 32'hed;
memory[390] = 32'hec;
memory[391] = 32'hf3;
memory[392] = 32'he4;
memory[393] = 32'hfa;
memory[394] = 32'hf9;
memory[395] = 32'hf8;
memory[396] = 32'hf7;
memory[397] = 32'hf6;
memory[398] = 32'hf5;
memory[399] = 32'hf4;
memory[400] = 32'hf3;
memory[401] = 32'hf2;
memory[402] = 32'hf1;
memory[403] = 32'hf0;
memory[404] = 32'hef;
memory[405] = 32'hee;
memory[406] = 32'hed;
memory[407] = 32'hec;
memory[408] = 32'heb;
memory[409] = 32'hea;
memory[410] = 32'he9;
memory[411] = 32'he8;
memory[412] = 32'he7;
memory[413] = 32'he6;
memory[414] = 32'he5;
memory[415] = 32'he4;
memory[416] = 32'he3;
memory[417] = 32'he2;
memory[418] = 32'he1;
memory[419] = 32'hfe;
memory[420] = 32'hfd;
memory[421] = 32'hfc;
memory[422] = 32'hfb;
memory[423] = 32'hfa;
memory[424] = 32'hf9;
memory[425] = 32'hf8;
memory[426] = 32'hf7;
memory[427] = 32'hf6;
memory[428] = 32'hf5;
memory[429] = 32'hf4;
memory[430] = 32'hf3;
memory[431] = 32'hf2;
memory[432] = 32'hf1;
memory[433] = 32'hf0;
memory[434] = 32'hef;
memory[435] = 32'hee;
memory[436] = 32'hed;
memory[437] = 32'hec;
memory[438] = 32'heb;
memory[439] = 32'hea;
memory[440] = 32'he9;
memory[441] = 32'he8;
memory[442] = 32'he7;
memory[443] = 32'he6;
memory[444] = 32'he5;
memory[445] = 32'he3;
memory[446] = 32'he6;
memory[447] = 32'hf1;
memory[448] = 32'he6;
memory[449] = 32'he3;
memory[450] = 32'he8;
memory[451] = 32'hf5;
memory[452] = 32'hf7;
memory[453] = 32'hee;
memory[454] = 32'hed;
memory[455] = 32'hf4;
memory[456] = 32'he5;
memory[457] = 32'hfc;
memory[458] = 32'hfc;
memory[459] = 32'hfb;
memory[460] = 32'hfa;
memory[461] = 32'hf9;
memory[462] = 32'hf8;
memory[463] = 32'hf7;
memory[464] = 32'hf6;
memory[465] = 32'hf5;
memory[466] = 32'hf4;
memory[467] = 32'hf3;
memory[468] = 32'hf2;
memory[469] = 32'hf1;
memory[470] = 32'hf0;
memory[471] = 32'hef;
memory[472] = 32'hee;
memory[473] = 32'hed;
memory[474] = 32'hec;
memory[475] = 32'heb;
memory[476] = 32'hea;
memory[477] = 32'he9;
memory[478] = 32'he8;
memory[479] = 32'he7;
memory[480] = 32'he6;
memory[481] = 32'he5;
memory[482] = 32'he4;
memory[483] = 32'he3;
memory[484] = 32'he2;
memory[485] = 32'he1;
memory[486] = 32'hfe;
memory[487] = 32'hfd;
memory[488] = 32'hfc;
memory[489] = 32'hfb;
memory[490] = 32'hfa;
memory[491] = 32'hf9;
memory[492] = 32'hf8;
memory[493] = 32'hf7;
memory[494] = 32'hf6;
memory[495] = 32'hf5;
memory[496] = 32'hf4;
memory[497] = 32'hf3;
memory[498] = 32'hf2;
memory[499] = 32'hf1;
memory[500] = 32'hf0;
memory[501] = 32'hef;
memory[502] = 32'hee;
memory[503] = 32'hed;
memory[504] = 32'hec;
memory[505] = 32'heb;
memory[506] = 32'hea;
memory[507] = 32'he9;
memory[508] = 32'he7;
memory[509] = 32'he2;
memory[510] = 32'he5;
memory[511] = 32'hf0;
memory[512] = 32'he5;
memory[513] = 32'he2;
memory[514] = 32'he7;
memory[515] = 32'hf4;
memory[516] = 32'hf8;
memory[517] = 32'hef;
memory[518] = 32'hee;
memory[519] = 32'hf5;
memory[520] = 32'he6;
memory[521] = 32'hfd;
memory[522] = 32'hfe;
memory[523] = 32'he8;
memory[524] = 32'he7;
memory[525] = 32'he6;
memory[526] = 32'he5;
memory[527] = 32'he4;
memory[528] = 32'he3;
memory[529] = 32'he2;
memory[530] = 32'he1;
memory[531] = 32'hfe;
memory[532] = 32'hfd;
memory[533] = 32'hfc;
memory[534] = 32'hfb;
memory[535] = 32'hfa;
memory[536] = 32'hf9;
memory[537] = 32'hf8;
memory[538] = 32'hf7;
memory[539] = 32'hf6;
memory[540] = 32'hf5;
memory[541] = 32'hf4;
memory[542] = 32'hf3;
memory[543] = 32'hf2;
memory[544] = 32'hf1;
memory[545] = 32'hf0;
memory[546] = 32'hef;
memory[547] = 32'hee;
memory[548] = 32'hed;
memory[549] = 32'hec;
memory[550] = 32'heb;
memory[551] = 32'hea;
memory[552] = 32'he9;
memory[553] = 32'he8;
memory[554] = 32'he7;
memory[555] = 32'he6;
memory[556] = 32'he5;
memory[557] = 32'he4;
memory[558] = 32'he3;
memory[559] = 32'he2;
memory[560] = 32'he1;
memory[561] = 32'hfe;
memory[562] = 32'hfd;
memory[563] = 32'hfc;
memory[564] = 32'hfb;
memory[565] = 32'hfa;
memory[566] = 32'hf9;
memory[567] = 32'hf8;
memory[568] = 32'hf7;
memory[569] = 32'hf6;
memory[570] = 32'hf5;
memory[571] = 32'hf3;
memory[572] = 32'he6;
memory[573] = 32'he1;
memory[574] = 32'he4;
memory[575] = 32'hef;
memory[576] = 32'he4;
memory[577] = 32'he1;
memory[578] = 32'he6;
memory[579] = 32'hf3;
memory[580] = 32'hf9;
memory[581] = 32'hf0;
memory[582] = 32'hef;
memory[583] = 32'hf6;
memory[584] = 32'he7;
memory[585] = 32'hfe;
memory[586] = 32'he1;
memory[587] = 32'hea;
memory[588] = 32'hfa;
memory[589] = 32'hf9;
memory[590] = 32'hf8;
memory[591] = 32'hf7;
memory[592] = 32'hf6;
memory[593] = 32'hf5;
memory[594] = 32'hf4;
memory[595] = 32'hf3;
memory[596] = 32'hf2;
memory[597] = 32'hf1;
memory[598] = 32'hf0;
memory[599] = 32'hef;
memory[600] = 32'hee;
memory[601] = 32'hed;
memory[602] = 32'hec;
memory[603] = 32'heb;
memory[604] = 32'hea;
memory[605] = 32'he9;
memory[606] = 32'he8;
memory[607] = 32'he7;
memory[608] = 32'he6;
memory[609] = 32'he5;
memory[610] = 32'he4;
memory[611] = 32'he3;
memory[612] = 32'he2;
memory[613] = 32'he1;
memory[614] = 32'hfe;
memory[615] = 32'hfd;
memory[616] = 32'hfc;
memory[617] = 32'hfb;
memory[618] = 32'hfa;
memory[619] = 32'hf9;
memory[620] = 32'hf8;
memory[621] = 32'hf7;
memory[622] = 32'hf6;
memory[623] = 32'hf5;
memory[624] = 32'hf4;
memory[625] = 32'hf3;
memory[626] = 32'hf2;
memory[627] = 32'hf1;
memory[628] = 32'hf0;
memory[629] = 32'hef;
memory[630] = 32'hee;
memory[631] = 32'hed;
memory[632] = 32'hec;
memory[633] = 32'heb;
memory[634] = 32'he9;
memory[635] = 32'hf2;
memory[636] = 32'he5;
memory[637] = 32'hfe;
memory[638] = 32'he3;
memory[639] = 32'hee;
memory[640] = 32'he3;
memory[641] = 32'hfe;
memory[642] = 32'he5;
memory[643] = 32'hf2;
memory[644] = 32'hfa;
memory[645] = 32'hf1;
memory[646] = 32'hf0;
memory[647] = 32'hf7;
memory[648] = 32'he8;
memory[649] = 32'he1;
memory[650] = 32'he2;
memory[651] = 32'heb;
memory[652] = 32'hfc;
memory[653] = 32'hf6;
memory[654] = 32'hf5;
memory[655] = 32'hf4;
memory[656] = 32'hf3;
memory[657] = 32'hf2;
memory[658] = 32'hf1;
memory[659] = 32'hf0;
memory[660] = 32'hef;
memory[661] = 32'hee;
memory[662] = 32'hed;
memory[663] = 32'hec;
memory[664] = 32'heb;
memory[665] = 32'hea;
memory[666] = 32'he9;
memory[667] = 32'he8;
memory[668] = 32'he7;
memory[669] = 32'he6;
memory[670] = 32'he5;
memory[671] = 32'he4;
memory[672] = 32'he3;
memory[673] = 32'he2;
memory[674] = 32'he1;
memory[675] = 32'hfe;
memory[676] = 32'hfd;
memory[677] = 32'hfc;
memory[678] = 32'hfb;
memory[679] = 32'hfa;
memory[680] = 32'hf9;
memory[681] = 32'hf8;
memory[682] = 32'hf7;
memory[683] = 32'hf6;
memory[684] = 32'hf5;
memory[685] = 32'hf4;
memory[686] = 32'hf3;
memory[687] = 32'hf2;
memory[688] = 32'hf1;
memory[689] = 32'hf0;
memory[690] = 32'hef;
memory[691] = 32'hee;
memory[692] = 32'hed;
memory[693] = 32'hec;
memory[694] = 32'heb;
memory[695] = 32'hea;
memory[696] = 32'he9;
memory[697] = 32'he7;
memory[698] = 32'he8;
memory[699] = 32'hf1;
memory[700] = 32'he4;
memory[701] = 32'hfd;
memory[702] = 32'he2;
memory[703] = 32'hed;
memory[704] = 32'he2;
memory[705] = 32'hfd;
memory[706] = 32'he4;
memory[707] = 32'hf1;
memory[708] = 32'hfb;
memory[709] = 32'hf2;
memory[710] = 32'hf1;
memory[711] = 32'hf8;
memory[712] = 32'he9;
memory[713] = 32'he2;
memory[714] = 32'he3;
memory[715] = 32'hec;
memory[716] = 32'hfd;
memory[717] = 32'hf8;
memory[718] = 32'hfa;
memory[719] = 32'hf9;
memory[720] = 32'hf8;
memory[721] = 32'hf7;
memory[722] = 32'hf6;
memory[723] = 32'hf5;
memory[724] = 32'hf4;
memory[725] = 32'hf3;
memory[726] = 32'hf2;
memory[727] = 32'hf1;
memory[728] = 32'hf0;
memory[729] = 32'hef;
memory[730] = 32'hee;
memory[731] = 32'hed;
memory[732] = 32'hec;
memory[733] = 32'heb;
memory[734] = 32'hea;
memory[735] = 32'he9;
memory[736] = 32'he8;
memory[737] = 32'he7;
memory[738] = 32'he6;
memory[739] = 32'he5;
memory[740] = 32'he4;
memory[741] = 32'he3;
memory[742] = 32'he2;
memory[743] = 32'he1;
memory[744] = 32'hfe;
memory[745] = 32'hfd;
memory[746] = 32'hfc;
memory[747] = 32'hfb;
memory[748] = 32'hfa;
memory[749] = 32'hf9;
memory[750] = 32'hf8;
memory[751] = 32'hf7;
memory[752] = 32'hf6;
memory[753] = 32'hf5;
memory[754] = 32'hf4;
memory[755] = 32'hf3;
memory[756] = 32'hf2;
memory[757] = 32'hf1;
memory[758] = 32'hf0;
memory[759] = 32'hef;
memory[760] = 32'hed;
memory[761] = 32'he6;
memory[762] = 32'he7;
memory[763] = 32'hf0;
memory[764] = 32'he3;
memory[765] = 32'hfc;
memory[766] = 32'he1;
memory[767] = 32'hec;
memory[768] = 32'he1;
memory[769] = 32'hfc;
memory[770] = 32'he3;
memory[771] = 32'hf0;
memory[772] = 32'hfc;
memory[773] = 32'hf3;
memory[774] = 32'hf2;
memory[775] = 32'hf9;
memory[776] = 32'hea;
memory[777] = 32'he3;
memory[778] = 32'he4;
memory[779] = 32'hed;
memory[780] = 32'hfe;
memory[781] = 32'hf9;
memory[782] = 32'hfc;
memory[783] = 32'he8;
memory[784] = 32'he7;
memory[785] = 32'he6;
memory[786] = 32'he5;
memory[787] = 32'he4;
memory[788] = 32'he3;
memory[789] = 32'he2;
memory[790] = 32'he1;
memory[791] = 32'hfe;
memory[792] = 32'hfd;
memory[793] = 32'hfc;
memory[794] = 32'hfb;
memory[795] = 32'hfa;
memory[796] = 32'hf9;
memory[797] = 32'hf8;
memory[798] = 32'hf7;
memory[799] = 32'hf6;
memory[800] = 32'hf5;
memory[801] = 32'hf4;
memory[802] = 32'hf3;
memory[803] = 32'hf2;
memory[804] = 32'hf1;
memory[805] = 32'hf0;
memory[806] = 32'hef;
memory[807] = 32'hee;
memory[808] = 32'hed;
memory[809] = 32'hec;
memory[810] = 32'heb;
memory[811] = 32'hea;
memory[812] = 32'he9;
memory[813] = 32'he8;
memory[814] = 32'he7;
memory[815] = 32'he6;
memory[816] = 32'he5;
memory[817] = 32'he4;
memory[818] = 32'he3;
memory[819] = 32'he2;
memory[820] = 32'he1;
memory[821] = 32'hfe;
memory[822] = 32'hfd;
memory[823] = 32'hfb;
memory[824] = 32'hec;
memory[825] = 32'he5;
memory[826] = 32'he6;
memory[827] = 32'hef;
memory[828] = 32'he2;
memory[829] = 32'hfb;
memory[830] = 32'hfe;
memory[831] = 32'heb;
memory[832] = 32'hfe;
memory[833] = 32'hfb;
memory[834] = 32'he2;
memory[835] = 32'hef;
memory[836] = 32'hfd;
memory[837] = 32'hf4;
memory[838] = 32'hf3;
memory[839] = 32'hfa;
memory[840] = 32'heb;
memory[841] = 32'he4;
memory[842] = 32'he5;
memory[843] = 32'hee;
memory[844] = 32'he1;
memory[845] = 32'hfa;
memory[846] = 32'hfd;
memory[847] = 32'hea;
memory[848] = 32'hfc;
memory[849] = 32'hfb;
memory[850] = 32'hfa;
memory[851] = 32'hf9;
memory[852] = 32'hf8;
memory[853] = 32'hf7;
memory[854] = 32'hf6;
memory[855] = 32'hf5;
memory[856] = 32'hf4;
memory[857] = 32'hf3;
memory[858] = 32'hf2;
memory[859] = 32'hf1;
memory[860] = 32'hf0;
memory[861] = 32'hef;
memory[862] = 32'hee;
memory[863] = 32'hed;
memory[864] = 32'hec;
memory[865] = 32'heb;
memory[866] = 32'hea;
memory[867] = 32'he9;
memory[868] = 32'he8;
memory[869] = 32'he7;
memory[870] = 32'he6;
memory[871] = 32'he5;
memory[872] = 32'he4;
memory[873] = 32'he3;
memory[874] = 32'he2;
memory[875] = 32'he1;
memory[876] = 32'hfe;
memory[877] = 32'hfd;
memory[878] = 32'hfc;
memory[879] = 32'hfb;
memory[880] = 32'hfa;
memory[881] = 32'hf9;
memory[882] = 32'hf8;
memory[883] = 32'hf7;
memory[884] = 32'hf6;
memory[885] = 32'hf5;
memory[886] = 32'hf3;
memory[887] = 32'hfa;
memory[888] = 32'heb;
memory[889] = 32'he4;
memory[890] = 32'he5;
memory[891] = 32'hee;
memory[892] = 32'he1;
memory[893] = 32'hfa;
memory[894] = 32'hfd;
memory[895] = 32'hea;
memory[896] = 32'hfd;
memory[897] = 32'hfa;
memory[898] = 32'he1;
memory[899] = 32'hee;
memory[900] = 32'hfe;
memory[901] = 32'hf5;
memory[902] = 32'hf4;
memory[903] = 32'hfb;
memory[904] = 32'hec;
memory[905] = 32'he5;
memory[906] = 32'he6;
memory[907] = 32'hef;
memory[908] = 32'he2;
memory[909] = 32'hfb;
memory[910] = 32'hfe;
memory[911] = 32'heb;
memory[912] = 32'hfe;
memory[913] = 32'hfa;
memory[914] = 32'hf9;
memory[915] = 32'hf8;
memory[916] = 32'hf7;
memory[917] = 32'hf6;
memory[918] = 32'hf5;
memory[919] = 32'hf4;
memory[920] = 32'hf3;
memory[921] = 32'hf2;
memory[922] = 32'hf1;
memory[923] = 32'hf0;
memory[924] = 32'hef;
memory[925] = 32'hee;
memory[926] = 32'hed;
memory[927] = 32'hec;
memory[928] = 32'heb;
memory[929] = 32'hea;
memory[930] = 32'he9;
memory[931] = 32'he8;
memory[932] = 32'he7;
memory[933] = 32'he6;
memory[934] = 32'he5;
memory[935] = 32'he4;
memory[936] = 32'he3;
memory[937] = 32'he2;
memory[938] = 32'he1;
memory[939] = 32'hfe;
memory[940] = 32'hfd;
memory[941] = 32'hfc;
memory[942] = 32'hfb;
memory[943] = 32'hfa;
memory[944] = 32'hf9;
memory[945] = 32'hf8;
memory[946] = 32'hf7;
memory[947] = 32'hf6;
memory[948] = 32'hf5;
memory[949] = 32'hf3;
memory[950] = 32'hf2;
memory[951] = 32'hf9;
memory[952] = 32'hea;
memory[953] = 32'he3;
memory[954] = 32'he4;
memory[955] = 32'hed;
memory[956] = 32'hfe;
memory[957] = 32'hf9;
memory[958] = 32'hfc;
memory[959] = 32'he9;
memory[960] = 32'hfc;
memory[961] = 32'hf9;
memory[962] = 32'hfe;
memory[963] = 32'hed;
memory[964] = 32'he1;
memory[965] = 32'hf6;
memory[966] = 32'hf5;
memory[967] = 32'hfc;
memory[968] = 32'hed;
memory[969] = 32'he6;
memory[970] = 32'he7;
memory[971] = 32'hf0;
memory[972] = 32'he3;
memory[973] = 32'hfc;
memory[974] = 32'he1;
memory[975] = 32'hec;
memory[976] = 32'he1;
memory[977] = 32'hfc;
memory[978] = 32'he2;
memory[979] = 32'he1;
memory[980] = 32'hfe;
memory[981] = 32'hfd;
memory[982] = 32'hfc;
memory[983] = 32'hfb;
memory[984] = 32'hfa;
memory[985] = 32'hf9;
memory[986] = 32'hf8;
memory[987] = 32'hf7;
memory[988] = 32'hf6;
memory[989] = 32'hf5;
memory[990] = 32'hf4;
memory[991] = 32'hf3;
memory[992] = 32'hf2;
memory[993] = 32'hf1;
memory[994] = 32'hf0;
memory[995] = 32'hef;
memory[996] = 32'hee;
memory[997] = 32'hed;
memory[998] = 32'hec;
memory[999] = 32'heb;
memory[1000] = 32'hea;
memory[1001] = 32'he9;
memory[1002] = 32'he8;
memory[1003] = 32'he7;
memory[1004] = 32'he6;
memory[1005] = 32'he5;
memory[1006] = 32'he4;
memory[1007] = 32'he3;
memory[1008] = 32'he2;
memory[1009] = 32'he1;
memory[1010] = 32'hfe;
memory[1011] = 32'hfd;
memory[1012] = 32'hfb;
memory[1013] = 32'hf2;
memory[1014] = 32'hf1;
memory[1015] = 32'hf8;
memory[1016] = 32'he9;
memory[1017] = 32'he2;
memory[1018] = 32'he3;
memory[1019] = 32'hec;
memory[1020] = 32'hfd;
memory[1021] = 32'hf8;
memory[1022] = 32'hfb;
memory[1023] = 32'he8;
memory[1024] = 32'hfb;
memory[1025] = 32'hf8;
memory[1026] = 32'hfd;
memory[1027] = 32'hec;
memory[1028] = 32'he2;
memory[1029] = 32'hf7;
memory[1030] = 32'hf6;
memory[1031] = 32'hfd;
memory[1032] = 32'hee;
memory[1033] = 32'he7;
memory[1034] = 32'he8;
memory[1035] = 32'hf1;
memory[1036] = 32'he4;
memory[1037] = 32'hfd;
memory[1038] = 32'he2;
memory[1039] = 32'hed;
memory[1040] = 32'he2;
memory[1041] = 32'hfd;
memory[1042] = 32'he4;
memory[1043] = 32'hf0;
memory[1044] = 32'hef;
memory[1045] = 32'hee;
memory[1046] = 32'hed;
memory[1047] = 32'hec;
memory[1048] = 32'heb;
memory[1049] = 32'hea;
memory[1050] = 32'he9;
memory[1051] = 32'he8;
memory[1052] = 32'he7;
memory[1053] = 32'he6;
memory[1054] = 32'he5;
memory[1055] = 32'he4;
memory[1056] = 32'he3;
memory[1057] = 32'he2;
memory[1058] = 32'he1;
memory[1059] = 32'hfe;
memory[1060] = 32'hfd;
memory[1061] = 32'hfc;
memory[1062] = 32'hfb;
memory[1063] = 32'hfa;
memory[1064] = 32'hf9;
memory[1065] = 32'hf8;
memory[1066] = 32'hf7;
memory[1067] = 32'hf6;
memory[1068] = 32'hf5;
memory[1069] = 32'hf4;
memory[1070] = 32'hf3;
memory[1071] = 32'hf2;
memory[1072] = 32'hf1;
memory[1073] = 32'hf0;
memory[1074] = 32'hef;
memory[1075] = 32'hed;
memory[1076] = 32'hfa;
memory[1077] = 32'hf1;
memory[1078] = 32'hf0;
memory[1079] = 32'hf7;
memory[1080] = 32'he8;
memory[1081] = 32'he1;
memory[1082] = 32'he2;
memory[1083] = 32'heb;
memory[1084] = 32'hfc;
memory[1085] = 32'hf7;
memory[1086] = 32'hfa;
memory[1087] = 32'he7;
memory[1088] = 32'hfa;
memory[1089] = 32'hf7;
memory[1090] = 32'hfc;
memory[1091] = 32'heb;
memory[1092] = 32'he3;
memory[1093] = 32'hf8;
memory[1094] = 32'hf7;
memory[1095] = 32'hfe;
memory[1096] = 32'hef;
memory[1097] = 32'he8;
memory[1098] = 32'he9;
memory[1099] = 32'hf2;
memory[1100] = 32'he5;
memory[1101] = 32'hfe;
memory[1102] = 32'he3;
memory[1103] = 32'hee;
memory[1104] = 32'he3;
memory[1105] = 32'hfe;
memory[1106] = 32'he5;
memory[1107] = 32'hf2;
memory[1108] = 32'he8;
memory[1109] = 32'he7;
memory[1110] = 32'he6;
memory[1111] = 32'he5;
memory[1112] = 32'he4;
memory[1113] = 32'he3;
memory[1114] = 32'he2;
memory[1115] = 32'he1;
memory[1116] = 32'hfe;
memory[1117] = 32'hfd;
memory[1118] = 32'hfc;
memory[1119] = 32'hfb;
memory[1120] = 32'hfa;
memory[1121] = 32'hf9;
memory[1122] = 32'hf8;
memory[1123] = 32'hf7;
memory[1124] = 32'hf6;
memory[1125] = 32'hf5;
memory[1126] = 32'hf4;
memory[1127] = 32'hf3;
memory[1128] = 32'hf2;
memory[1129] = 32'hf1;
memory[1130] = 32'hf0;
memory[1131] = 32'hef;
memory[1132] = 32'hee;
memory[1133] = 32'hed;
memory[1134] = 32'hec;
memory[1135] = 32'heb;
memory[1136] = 32'hea;
memory[1137] = 32'he9;
memory[1138] = 32'he7;
memory[1139] = 32'hec;
memory[1140] = 32'hf9;
memory[1141] = 32'hf0;
memory[1142] = 32'hef;
memory[1143] = 32'hf6;
memory[1144] = 32'he7;
memory[1145] = 32'hfe;
memory[1146] = 32'he1;
memory[1147] = 32'hea;
memory[1148] = 32'hfb;
memory[1149] = 32'hf6;
memory[1150] = 32'hf9;
memory[1151] = 32'he6;
memory[1152] = 32'hf9;
memory[1153] = 32'hf6;
memory[1154] = 32'hfb;
memory[1155] = 32'hea;
memory[1156] = 32'he4;
memory[1157] = 32'hf9;
memory[1158] = 32'hf8;
memory[1159] = 32'he1;
memory[1160] = 32'hf0;
memory[1161] = 32'he9;
memory[1162] = 32'hea;
memory[1163] = 32'hf3;
memory[1164] = 32'he6;
memory[1165] = 32'he1;
memory[1166] = 32'he4;
memory[1167] = 32'hef;
memory[1168] = 32'he4;
memory[1169] = 32'he1;
memory[1170] = 32'he6;
memory[1171] = 32'hf3;
memory[1172] = 32'hea;
memory[1173] = 32'he8;
memory[1174] = 32'he7;
memory[1175] = 32'he6;
memory[1176] = 32'he5;
memory[1177] = 32'he4;
memory[1178] = 32'he3;
memory[1179] = 32'he2;
memory[1180] = 32'he1;
memory[1181] = 32'hfe;
memory[1182] = 32'hfd;
memory[1183] = 32'hfc;
memory[1184] = 32'hfb;
memory[1185] = 32'hfa;
memory[1186] = 32'hf9;
memory[1187] = 32'hf8;
memory[1188] = 32'hf7;
memory[1189] = 32'hf6;
memory[1190] = 32'hf5;
memory[1191] = 32'hf4;
memory[1192] = 32'hf3;
memory[1193] = 32'hf2;
memory[1194] = 32'hf1;
memory[1195] = 32'hf0;
memory[1196] = 32'hef;
memory[1197] = 32'hee;
memory[1198] = 32'hed;
memory[1199] = 32'hec;
memory[1200] = 32'heb;
memory[1201] = 32'he9;
memory[1202] = 32'he6;
memory[1203] = 32'heb;
memory[1204] = 32'hf8;
memory[1205] = 32'hef;
memory[1206] = 32'hee;
memory[1207] = 32'hf5;
memory[1208] = 32'he6;
memory[1209] = 32'hfd;
memory[1210] = 32'hfe;
memory[1211] = 32'he9;
memory[1212] = 32'hfa;
memory[1213] = 32'hf5;
memory[1214] = 32'hf8;
memory[1215] = 32'he5;
memory[1216] = 32'hf8;
memory[1217] = 32'hf5;
memory[1218] = 32'hfa;
memory[1219] = 32'he9;
memory[1220] = 32'he5;
memory[1221] = 32'hfa;
memory[1222] = 32'hf9;
memory[1223] = 32'he2;
memory[1224] = 32'hf1;
memory[1225] = 32'hea;
memory[1226] = 32'heb;
memory[1227] = 32'hf4;
memory[1228] = 32'he7;
memory[1229] = 32'he2;
memory[1230] = 32'he5;
memory[1231] = 32'hf0;
memory[1232] = 32'he5;
memory[1233] = 32'he2;
memory[1234] = 32'he7;
memory[1235] = 32'hf4;
memory[1236] = 32'heb;
memory[1237] = 32'hea;
memory[1238] = 32'hf0;
memory[1239] = 32'h65;
memory[1240] = 32'h65;
memory[1241] = 32'h65;
memory[1242] = 32'h65;
memory[1243] = 32'heb;
memory[1244] = 32'hea;
memory[1245] = 32'he9;
memory[1246] = 32'he8;
memory[1247] = 32'he7;
memory[1248] = 32'he6;
memory[1249] = 32'he5;
memory[1250] = 32'he4;
memory[1251] = 32'he3;
memory[1252] = 32'he2;
memory[1253] = 32'he1;
memory[1254] = 32'hfe;
memory[1255] = 32'hfd;
memory[1256] = 32'hfc;
memory[1257] = 32'hfb;
memory[1258] = 32'hfa;
memory[1259] = 32'hf9;
memory[1260] = 32'hf8;
memory[1261] = 32'hf7;
memory[1262] = 32'hf6;
memory[1263] = 32'hf5;
memory[1264] = 32'hf3;
memory[1265] = 32'he8;
memory[1266] = 32'he5;
memory[1267] = 32'hea;
memory[1268] = 32'hf7;
memory[1269] = 32'hee;
memory[1270] = 32'hed;
memory[1271] = 32'hf4;
memory[1272] = 32'he5;
memory[1273] = 32'hfc;
memory[1274] = 32'hfd;
memory[1275] = 32'he8;
memory[1276] = 32'hf9;
memory[1277] = 32'hf4;
memory[1278] = 32'hf7;
memory[1279] = 32'he4;
memory[1280] = 32'hf7;
memory[1281] = 32'hf4;
memory[1282] = 32'hf9;
memory[1283] = 32'he8;
memory[1284] = 32'he6;
memory[1285] = 32'hfb;
memory[1286] = 32'hfa;
memory[1287] = 32'he3;
memory[1288] = 32'hf2;
memory[1289] = 32'heb;
memory[1290] = 32'hec;
memory[1291] = 32'hf5;
memory[1292] = 32'he8;
memory[1293] = 32'he3;
memory[1294] = 32'he6;
memory[1295] = 32'hf1;
memory[1296] = 32'he6;
memory[1297] = 32'he3;
memory[1298] = 32'he8;
memory[1299] = 32'hf5;
memory[1300] = 32'hec;
memory[1301] = 32'heb;
memory[1302] = 32'hf2;
memory[1303] = 32'h65;
memory[1304] = 32'h65;
memory[1305] = 32'h65;
memory[1306] = 32'h65;
memory[1307] = 32'hfc;
memory[1308] = 32'hfb;
memory[1309] = 32'hfa;
memory[1310] = 32'hf9;
memory[1311] = 32'hf8;
memory[1312] = 32'hf7;
memory[1313] = 32'hf6;
memory[1314] = 32'hf5;
memory[1315] = 32'hf4;
memory[1316] = 32'hf3;
memory[1317] = 32'hf2;
memory[1318] = 32'hf1;
memory[1319] = 32'hf0;
memory[1320] = 32'hef;
memory[1321] = 32'hee;
memory[1322] = 32'hed;
memory[1323] = 32'hec;
memory[1324] = 32'heb;
memory[1325] = 32'hea;
memory[1326] = 32'he9;
memory[1327] = 32'he7;
memory[1328] = 32'hf2;
memory[1329] = 32'he7;
memory[1330] = 32'he4;
memory[1331] = 32'he9;
memory[1332] = 32'hf6;
memory[1333] = 32'hed;
memory[1334] = 32'hec;
memory[1335] = 32'hf3;
memory[1336] = 32'he4;
memory[1337] = 32'hfb;
memory[1338] = 32'hfc;
memory[1339] = 32'he7;
memory[1340] = 32'hf8;
memory[1341] = 32'hf3;
memory[1342] = 32'hf6;
memory[1343] = 32'he3;
memory[1344] = 32'hf6;
memory[1345] = 32'hf3;
memory[1346] = 32'hf8;
memory[1347] = 32'he7;
memory[1348] = 32'he7;
memory[1349] = 32'hfc;
memory[1350] = 32'hfb;
memory[1351] = 32'he4;
memory[1352] = 32'hf3;
memory[1353] = 32'hec;
memory[1354] = 32'hed;
memory[1355] = 32'hf6;
memory[1356] = 32'he9;
memory[1357] = 32'he4;
memory[1358] = 32'he7;
memory[1359] = 32'hf2;
memory[1360] = 32'he7;
memory[1361] = 32'he4;
memory[1362] = 32'he9;
memory[1363] = 32'hf6;
memory[1364] = 32'hed;
memory[1365] = 32'hec;
memory[1366] = 32'hf3;
memory[1367] = 32'h65;
memory[1368] = 32'h65;
memory[1369] = 32'h65;
memory[1370] = 32'h65;
memory[1371] = 32'hf7;
memory[1372] = 32'hf6;
memory[1373] = 32'hf5;
memory[1374] = 32'hf4;
memory[1375] = 32'hf3;
memory[1376] = 32'hf2;
memory[1377] = 32'hf1;
memory[1378] = 32'hf0;
memory[1379] = 32'hef;
memory[1380] = 32'hee;
memory[1381] = 32'hed;
memory[1382] = 32'hec;
memory[1383] = 32'heb;
memory[1384] = 32'hea;
memory[1385] = 32'he9;
memory[1386] = 32'he8;
memory[1387] = 32'he7;
memory[1388] = 32'he6;
memory[1389] = 32'he5;
memory[1390] = 32'he3;
memory[1391] = 32'he6;
memory[1392] = 32'hf1;
memory[1393] = 32'he6;
memory[1394] = 32'he3;
memory[1395] = 32'he8;
memory[1396] = 32'hf5;
memory[1397] = 32'hec;
memory[1398] = 32'heb;
memory[1399] = 32'hf2;
memory[1400] = 32'he3;
memory[1401] = 32'hfa;
memory[1402] = 32'hfb;
memory[1403] = 32'he6;
memory[1404] = 32'hf7;
memory[1405] = 32'hf2;
memory[1406] = 32'hf5;
memory[1407] = 32'he2;
memory[1408] = 32'hf5;
memory[1409] = 32'hf2;
memory[1410] = 32'hf7;
memory[1411] = 32'he6;
memory[1412] = 32'he8;
memory[1413] = 32'hfd;
memory[1414] = 32'hfc;
memory[1415] = 32'he5;
memory[1416] = 32'hf4;
memory[1417] = 32'hed;
memory[1418] = 32'hee;
memory[1419] = 32'hf7;
memory[1420] = 32'hea;
memory[1421] = 32'he5;
memory[1422] = 32'he8;
memory[1423] = 32'hf3;
memory[1424] = 32'he8;
memory[1425] = 32'he5;
memory[1426] = 32'hea;
memory[1427] = 32'hf7;
memory[1428] = 32'hee;
memory[1429] = 32'hed;
memory[1430] = 32'hf4;
memory[1431] = 32'h65;
memory[1432] = 32'h65;
memory[1433] = 32'h65;
memory[1434] = 32'h65;
memory[1435] = 32'hfa;
memory[1436] = 32'hf9;
memory[1437] = 32'hf8;
memory[1438] = 32'hf7;
memory[1439] = 32'hf6;
memory[1440] = 32'hf5;
memory[1441] = 32'hf4;
memory[1442] = 32'hf3;
memory[1443] = 32'hf2;
memory[1444] = 32'hf1;
memory[1445] = 32'hf0;
memory[1446] = 32'hef;
memory[1447] = 32'hee;
memory[1448] = 32'hed;
memory[1449] = 32'hec;
memory[1450] = 32'heb;
memory[1451] = 32'hea;
memory[1452] = 32'he9;
memory[1453] = 32'he7;
memory[1454] = 32'he2;
memory[1455] = 32'he5;
memory[1456] = 32'hf0;
memory[1457] = 32'he5;
memory[1458] = 32'he2;
memory[1459] = 32'he7;
memory[1460] = 32'hf4;
memory[1461] = 32'heb;
memory[1462] = 32'hea;
memory[1463] = 32'hf1;
memory[1464] = 32'he2;
memory[1465] = 32'hf9;
memory[1466] = 32'hfa;
memory[1467] = 32'he5;
memory[1468] = 32'hf6;
memory[1469] = 32'hf1;
memory[1470] = 32'hf4;
memory[1471] = 32'he1;
memory[1472] = 32'hf4;
memory[1473] = 32'hf1;
memory[1474] = 32'hf6;
memory[1475] = 32'he5;
memory[1476] = 32'he9;
memory[1477] = 32'hfe;
memory[1478] = 32'hfd;
memory[1479] = 32'he6;
memory[1480] = 32'hf5;
memory[1481] = 32'hee;
memory[1482] = 32'hef;
memory[1483] = 32'hf8;
memory[1484] = 32'heb;
memory[1485] = 32'he6;
memory[1486] = 32'he9;
memory[1487] = 32'hf4;
memory[1488] = 32'he9;
memory[1489] = 32'he6;
memory[1490] = 32'heb;
memory[1491] = 32'hf8;
memory[1492] = 32'hef;
memory[1493] = 32'hee;
memory[1494] = 32'hf5;
memory[1495] = 32'he6;
memory[1496] = 32'hfd;
memory[1497] = 32'hfe;
memory[1498] = 32'he8;
memory[1499] = 32'he7;
memory[1500] = 32'he6;
memory[1501] = 32'he5;
memory[1502] = 32'he4;
memory[1503] = 32'he3;
memory[1504] = 32'he2;
memory[1505] = 32'he1;
memory[1506] = 32'hfe;
memory[1507] = 32'hfd;
memory[1508] = 32'hfc;
memory[1509] = 32'hfb;
memory[1510] = 32'hfa;
memory[1511] = 32'hf9;
memory[1512] = 32'hf8;
memory[1513] = 32'hf7;
memory[1514] = 32'hf6;
memory[1515] = 32'hf5;
memory[1516] = 32'hf3;
memory[1517] = 32'he6;
memory[1518] = 32'he1;
memory[1519] = 32'he4;
memory[1520] = 32'hef;
memory[1521] = 32'he4;
memory[1522] = 32'he1;
memory[1523] = 32'he6;
memory[1524] = 32'hf3;
memory[1525] = 32'hea;
memory[1526] = 32'he9;
memory[1527] = 32'hf0;
memory[1528] = 32'he1;
memory[1529] = 32'hf8;
memory[1530] = 32'hf9;
memory[1531] = 32'he4;
memory[1532] = 32'hf5;
memory[1533] = 32'hf0;
memory[1534] = 32'hf3;
memory[1535] = 32'hfe;
memory[1536] = 32'hf3;
memory[1537] = 32'hf0;
memory[1538] = 32'hf5;
memory[1539] = 32'he4;
memory[1540] = 32'hea;
memory[1541] = 32'he1;
memory[1542] = 32'hfe;
memory[1543] = 32'he7;
memory[1544] = 32'hf6;
memory[1545] = 32'hef;
memory[1546] = 32'hf0;
memory[1547] = 32'hf9;
memory[1548] = 32'hec;
memory[1549] = 32'he7;
memory[1550] = 32'hea;
memory[1551] = 32'hf5;
memory[1552] = 32'hea;
memory[1553] = 32'he7;
memory[1554] = 32'hec;
memory[1555] = 32'hf9;
memory[1556] = 32'hf0;
memory[1557] = 32'hef;
memory[1558] = 32'hf6;
memory[1559] = 32'he7;
memory[1560] = 32'hfe;
memory[1561] = 32'he1;
memory[1562] = 32'hea;
memory[1563] = 32'hfa;
memory[1564] = 32'hf9;
memory[1565] = 32'hf8;
memory[1566] = 32'hf7;
memory[1567] = 32'hf6;
memory[1568] = 32'hf5;
memory[1569] = 32'hf4;
memory[1570] = 32'hf3;
memory[1571] = 32'hf2;
memory[1572] = 32'hf1;
memory[1573] = 32'hf0;
memory[1574] = 32'hef;
memory[1575] = 32'hee;
memory[1576] = 32'hed;
memory[1577] = 32'hec;
memory[1578] = 32'heb;
memory[1579] = 32'he9;
memory[1580] = 32'hf2;
memory[1581] = 32'he5;
memory[1582] = 32'hfe;
memory[1583] = 32'he3;
memory[1584] = 32'hee;
memory[1585] = 32'he3;
memory[1586] = 32'hfe;
memory[1587] = 32'he5;
memory[1588] = 32'hf2;
memory[1589] = 32'he9;
memory[1590] = 32'he8;
memory[1591] = 32'hef;
memory[1592] = 32'hfe;
memory[1593] = 32'hf7;
memory[1594] = 32'hf8;
memory[1595] = 32'he3;
memory[1596] = 32'hf4;
memory[1597] = 32'hef;
memory[1598] = 32'hf2;
memory[1599] = 32'hfd;
memory[1600] = 32'hf2;
memory[1601] = 32'hef;
memory[1602] = 32'hf4;
memory[1603] = 32'he3;
memory[1604] = 32'heb;
memory[1605] = 32'he2;
memory[1606] = 32'he1;
memory[1607] = 32'he8;
memory[1608] = 32'hf7;
memory[1609] = 32'hf0;
memory[1610] = 32'hf1;
memory[1611] = 32'hfa;
memory[1612] = 32'hed;
memory[1613] = 32'he8;
memory[1614] = 32'heb;
memory[1615] = 32'hf6;
memory[1616] = 32'heb;
memory[1617] = 32'he8;
memory[1618] = 32'hed;
memory[1619] = 32'hfa;
memory[1620] = 32'hf1;
memory[1621] = 32'hf0;
memory[1622] = 32'hf7;
memory[1623] = 32'he8;
memory[1624] = 32'he1;
memory[1625] = 32'he2;
memory[1626] = 32'heb;
memory[1627] = 32'hfc;
memory[1628] = 32'hf6;
memory[1629] = 32'hf5;
memory[1630] = 32'hf4;
memory[1631] = 32'hf3;
memory[1632] = 32'hf2;
memory[1633] = 32'hf1;
memory[1634] = 32'hf0;
memory[1635] = 32'hef;
memory[1636] = 32'hee;
memory[1637] = 32'hed;
memory[1638] = 32'hec;
memory[1639] = 32'heb;
memory[1640] = 32'hea;
memory[1641] = 32'he9;
memory[1642] = 32'he7;
memory[1643] = 32'he8;
memory[1644] = 32'hf1;
memory[1645] = 32'he4;
memory[1646] = 32'hfd;
memory[1647] = 32'he2;
memory[1648] = 32'hed;
memory[1649] = 32'he2;
memory[1650] = 32'hfd;
memory[1651] = 32'he4;
memory[1652] = 32'hf1;
memory[1653] = 32'he8;
memory[1654] = 32'he7;
memory[1655] = 32'hee;
memory[1656] = 32'hfd;
memory[1657] = 32'hf6;
memory[1658] = 32'hf7;
memory[1659] = 32'he2;
memory[1660] = 32'hf3;
memory[1661] = 32'hee;
memory[1662] = 32'hf1;
memory[1663] = 32'hfc;
memory[1664] = 32'hf1;
memory[1665] = 32'hee;
memory[1666] = 32'hf3;
memory[1667] = 32'he2;
memory[1668] = 32'hec;
memory[1669] = 32'he3;
memory[1670] = 32'he2;
memory[1671] = 32'he9;
memory[1672] = 32'hf8;
memory[1673] = 32'hf1;
memory[1674] = 32'hf2;
memory[1675] = 32'hfb;
memory[1676] = 32'hee;
memory[1677] = 32'he9;
memory[1678] = 32'hec;
memory[1679] = 32'hf7;
memory[1680] = 32'hec;
memory[1681] = 32'he9;
memory[1682] = 32'hee;
memory[1683] = 32'hfb;
memory[1684] = 32'hf2;
memory[1685] = 32'hf1;
memory[1686] = 32'hf8;
memory[1687] = 32'he9;
memory[1688] = 32'he2;
memory[1689] = 32'he3;
memory[1690] = 32'hec;
memory[1691] = 32'hfd;
memory[1692] = 32'hf8;
memory[1693] = 32'hfa;
memory[1694] = 32'hf9;
memory[1695] = 32'hf8;
memory[1696] = 32'hf7;
memory[1697] = 32'hf6;
memory[1698] = 32'hf5;
memory[1699] = 32'hf4;
memory[1700] = 32'hf3;
memory[1701] = 32'hf2;
memory[1702] = 32'hf1;
memory[1703] = 32'hf0;
memory[1704] = 32'hef;
memory[1705] = 32'hed;
memory[1706] = 32'he6;
memory[1707] = 32'he7;
memory[1708] = 32'hf0;
memory[1709] = 32'he3;
memory[1710] = 32'hfc;
memory[1711] = 32'he1;
memory[1712] = 32'hec;
memory[1713] = 32'he1;
memory[1714] = 32'hfc;
memory[1715] = 32'he3;
memory[1716] = 32'hf0;
memory[1717] = 32'he7;
memory[1718] = 32'he6;
memory[1719] = 32'hed;
memory[1720] = 32'hfc;
memory[1721] = 32'hf5;
memory[1722] = 32'hf6;
memory[1723] = 32'he1;
memory[1724] = 32'hf2;
memory[1725] = 32'hed;
memory[1726] = 32'hf0;
memory[1727] = 32'hfb;
memory[1728] = 32'hf0;
memory[1729] = 32'hed;
memory[1730] = 32'hf2;
memory[1731] = 32'he1;
memory[1732] = 32'hed;
memory[1733] = 32'he4;
memory[1734] = 32'he3;
memory[1735] = 32'hea;
memory[1736] = 32'hf9;
memory[1737] = 32'hf2;
memory[1738] = 32'hf3;
memory[1739] = 32'hfc;
memory[1740] = 32'hef;
memory[1741] = 32'hea;
memory[1742] = 32'hed;
memory[1743] = 32'hf8;
memory[1744] = 32'hed;
memory[1745] = 32'hea;
memory[1746] = 32'hef;
memory[1747] = 32'hfc;
memory[1748] = 32'hf3;
memory[1749] = 32'hf2;
memory[1750] = 32'hf9;
memory[1751] = 32'hea;
memory[1752] = 32'he3;
memory[1753] = 32'he4;
memory[1754] = 32'hed;
memory[1755] = 32'hfe;
memory[1756] = 32'hf9;
memory[1757] = 32'hfc;
memory[1758] = 32'he8;
memory[1759] = 32'he7;
memory[1760] = 32'he6;
memory[1761] = 32'he5;
memory[1762] = 32'he4;
memory[1763] = 32'he3;
memory[1764] = 32'he2;
memory[1765] = 32'he1;
memory[1766] = 32'h64;
memory[1767] = 32'h64;
memory[1768] = 32'h64;
memory[1769] = 32'h64;
memory[1770] = 32'he5;
memory[1771] = 32'he6;
memory[1772] = 32'hef;
memory[1773] = 32'he2;
memory[1774] = 32'hfb;
memory[1775] = 32'hfe;
memory[1776] = 32'heb;
memory[1777] = 32'hfe;
memory[1778] = 32'hfb;
memory[1779] = 32'he2;
memory[1780] = 32'hef;
memory[1781] = 32'he6;
memory[1782] = 32'he5;
memory[1783] = 32'hec;
memory[1784] = 32'hfb;
memory[1785] = 32'hf4;
memory[1786] = 32'hf5;
memory[1787] = 32'hfe;
memory[1788] = 32'hf1;
memory[1789] = 32'hec;
memory[1790] = 32'hef;
memory[1791] = 32'hfa;
memory[1792] = 32'hef;
memory[1793] = 32'hec;
memory[1794] = 32'hf1;
memory[1795] = 32'hfe;
memory[1796] = 32'hee;
memory[1797] = 32'he5;
memory[1798] = 32'he4;
memory[1799] = 32'heb;
memory[1800] = 32'hfa;
memory[1801] = 32'hf3;
memory[1802] = 32'hf4;
memory[1803] = 32'hfd;
memory[1804] = 32'hf0;
memory[1805] = 32'heb;
memory[1806] = 32'hee;
memory[1807] = 32'hf9;
memory[1808] = 32'hee;
memory[1809] = 32'heb;
memory[1810] = 32'hf0;
memory[1811] = 32'hfd;
memory[1812] = 32'hf4;
memory[1813] = 32'hf3;
memory[1814] = 32'hfa;
memory[1815] = 32'heb;
memory[1816] = 32'he4;
memory[1817] = 32'he5;
memory[1818] = 32'hee;
memory[1819] = 32'he1;
memory[1820] = 32'hfa;
memory[1821] = 32'hfd;
memory[1822] = 32'hea;
memory[1823] = 32'hfc;
memory[1824] = 32'hfb;
memory[1825] = 32'hfa;
memory[1826] = 32'hf9;
memory[1827] = 32'hf8;
memory[1828] = 32'hf7;
memory[1829] = 32'hf6;
memory[1830] = 32'h64;
memory[1831] = 32'h63;
memory[1832] = 32'h64;
memory[1833] = 32'h64;
memory[1834] = 32'he4;
memory[1835] = 32'he5;
memory[1836] = 32'hee;
memory[1837] = 32'he1;
memory[1838] = 32'hfa;
memory[1839] = 32'hfd;
memory[1840] = 32'hea;
memory[1841] = 32'hfd;
memory[1842] = 32'hfa;
memory[1843] = 32'he1;
memory[1844] = 32'hee;
memory[1845] = 32'he5;
memory[1846] = 32'he4;
memory[1847] = 32'heb;
memory[1848] = 32'hfa;
memory[1849] = 32'hf3;
memory[1850] = 32'hf4;
memory[1851] = 32'hfd;
memory[1852] = 32'hf0;
memory[1853] = 32'heb;
memory[1854] = 32'hee;
memory[1855] = 32'hf9;
memory[1856] = 32'hee;
memory[1857] = 32'heb;
memory[1858] = 32'hf0;
memory[1859] = 32'hfd;
memory[1860] = 32'hef;
memory[1861] = 32'he6;
memory[1862] = 32'he5;
memory[1863] = 32'hec;
memory[1864] = 32'hfb;
memory[1865] = 32'hf4;
memory[1866] = 32'hf5;
memory[1867] = 32'hfe;
memory[1868] = 32'hf1;
memory[1869] = 32'hec;
memory[1870] = 32'hef;
memory[1871] = 32'hfa;
memory[1872] = 32'hef;
memory[1873] = 32'hec;
memory[1874] = 32'hf1;
memory[1875] = 32'hfe;
memory[1876] = 32'hf5;
memory[1877] = 32'hf4;
memory[1878] = 32'hfb;
memory[1879] = 32'hec;
memory[1880] = 32'he5;
memory[1881] = 32'he6;
memory[1882] = 32'hef;
memory[1883] = 32'he2;
memory[1884] = 32'hfb;
memory[1885] = 32'hfe;
memory[1886] = 32'heb;
memory[1887] = 32'hfe;
memory[1888] = 32'hfa;
memory[1889] = 32'hf9;
memory[1890] = 32'hf8;
memory[1891] = 32'h78;
memory[1892] = 32'h78;
memory[1893] = 32'hf5;
memory[1894] = 32'h64;
memory[1895] = 32'h64;
memory[1896] = 32'h63;
memory[1897] = 32'h64;
memory[1898] = 32'he3;
memory[1899] = 32'he4;
memory[1900] = 32'hed;
memory[1901] = 32'hfe;
memory[1902] = 32'hf9;
memory[1903] = 32'hfc;
memory[1904] = 32'he9;
memory[1905] = 32'hfc;
memory[1906] = 32'hf9;
memory[1907] = 32'hfe;
memory[1908] = 32'hed;
memory[1909] = 32'he4;
memory[1910] = 32'he3;
memory[1911] = 32'hea;
memory[1912] = 32'hf9;
memory[1913] = 32'hf2;
memory[1914] = 32'hf3;
memory[1915] = 32'hfc;
memory[1916] = 32'hef;
memory[1917] = 32'hea;
memory[1918] = 32'hed;
memory[1919] = 32'hf8;
memory[1920] = 32'hed;
memory[1921] = 32'hea;
memory[1922] = 32'hef;
memory[1923] = 32'hfc;
memory[1924] = 32'hf0;
memory[1925] = 32'he7;
memory[1926] = 32'he6;
memory[1927] = 32'hed;
memory[1928] = 32'hfc;
memory[1929] = 32'hf5;
memory[1930] = 32'hf6;
memory[1931] = 32'he1;
memory[1932] = 32'hf2;
memory[1933] = 32'hed;
memory[1934] = 32'hf0;
memory[1935] = 32'hfb;
memory[1936] = 32'hf0;
memory[1937] = 32'hed;
memory[1938] = 32'hf2;
memory[1939] = 32'he1;
memory[1940] = 32'hf6;
memory[1941] = 32'hf5;
memory[1942] = 32'hfc;
memory[1943] = 32'hed;
memory[1944] = 32'he6;
memory[1945] = 32'he7;
memory[1946] = 32'hf0;
memory[1947] = 32'he3;
memory[1948] = 32'hfc;
memory[1949] = 32'he1;
memory[1950] = 32'hec;
memory[1951] = 32'he1;
memory[1952] = 32'hfc;
memory[1953] = 32'he2;
memory[1954] = 32'he1;
memory[1955] = 32'h78;
memory[1956] = 32'h78;
memory[1957] = 32'h78;
memory[1958] = 32'h64;
memory[1959] = 32'h64;
memory[1960] = 32'h64;
memory[1961] = 32'h64;
memory[1962] = 32'he2;
memory[1963] = 32'he3;
memory[1964] = 32'hec;
memory[1965] = 32'hfd;
memory[1966] = 32'hf8;
memory[1967] = 32'hfb;
memory[1968] = 32'he8;
memory[1969] = 32'hfb;
memory[1970] = 32'hf8;
memory[1971] = 32'hfd;
memory[1972] = 32'hec;
memory[1973] = 32'he3;
memory[1974] = 32'he2;
memory[1975] = 32'he9;
memory[1976] = 32'hf8;
memory[1977] = 32'hf1;
memory[1978] = 32'hf2;
memory[1979] = 32'hfb;
memory[1980] = 32'hee;
memory[1981] = 32'he9;
memory[1982] = 32'hec;
memory[1983] = 32'hf7;
memory[1984] = 32'hec;
memory[1985] = 32'he9;
memory[1986] = 32'hee;
memory[1987] = 32'hfb;
memory[1988] = 32'hf1;
memory[1989] = 32'he8;
memory[1990] = 32'he7;
memory[1991] = 32'hee;
memory[1992] = 32'hfd;
memory[1993] = 32'hf6;
memory[1994] = 32'hf7;
memory[1995] = 32'he2;
memory[1996] = 32'hf3;
memory[1997] = 32'hee;
memory[1998] = 32'hf1;
memory[1999] = 32'hfc;
memory[2000] = 32'hf1;
memory[2001] = 32'hee;
memory[2002] = 32'hf3;
memory[2003] = 32'he2;
memory[2004] = 32'hf7;
memory[2005] = 32'hf6;
memory[2006] = 32'hfd;
memory[2007] = 32'hee;
memory[2008] = 32'he7;
memory[2009] = 32'he8;
memory[2010] = 32'hf1;
memory[2011] = 32'he4;
memory[2012] = 32'hfd;
memory[2013] = 32'he2;
memory[2014] = 32'hed;
memory[2015] = 32'he2;
memory[2016] = 32'hfd;
memory[2017] = 32'he4;
memory[2018] = 32'hf0;
memory[2019] = 32'hef;
memory[2020] = 32'hed;
memory[2021] = 32'hfa;
memory[2022] = 32'hf1;
memory[2023] = 32'hf0;
memory[2024] = 32'hf7;
memory[2025] = 32'he8;
memory[2026] = 32'he1;
memory[2027] = 32'he2;
memory[2028] = 32'heb;
memory[2029] = 32'hfc;
memory[2030] = 32'hf7;
memory[2031] = 32'hfa;
memory[2032] = 32'he7;
memory[2033] = 32'hfa;
memory[2034] = 32'hf7;
memory[2035] = 32'hfc;
memory[2036] = 32'heb;
memory[2037] = 32'he2;
memory[2038] = 32'he1;
memory[2039] = 32'he8;
memory[2040] = 32'hf7;
memory[2041] = 32'hf0;
memory[2042] = 32'hf1;
memory[2043] = 32'hfa;
memory[2044] = 32'hed;
memory[2045] = 32'he8;
memory[2046] = 32'heb;
memory[2047] = 32'hf6;
memory[2048] = 32'heb;
memory[2049] = 32'he8;
memory[2050] = 32'hed;
memory[2051] = 32'hfa;
memory[2052] = 32'hf2;
memory[2053] = 32'he9;
memory[2054] = 32'he8;
memory[2055] = 32'hef;
memory[2056] = 32'hfe;
memory[2057] = 32'hf7;
memory[2058] = 32'hf8;
memory[2059] = 32'he3;
memory[2060] = 32'hf4;
memory[2061] = 32'hef;
memory[2062] = 32'hf2;
memory[2063] = 32'hfd;
memory[2064] = 32'hf2;
memory[2065] = 32'hef;
memory[2066] = 32'hf4;
memory[2067] = 32'he3;
memory[2068] = 32'hf8;
memory[2069] = 32'hf7;
memory[2070] = 32'hfe;
memory[2071] = 32'hef;
memory[2072] = 32'he8;
memory[2073] = 32'he9;
memory[2074] = 32'hf2;
memory[2075] = 32'he5;
memory[2076] = 32'hfe;
memory[2077] = 32'he3;
memory[2078] = 32'hee;
memory[2079] = 32'he3;
memory[2080] = 32'hfe;
memory[2081] = 32'he5;
memory[2082] = 32'h65;
memory[2083] = 32'h78;
memory[2084] = 32'h78;
memory[2085] = 32'h78;
memory[2086] = 32'h78;
memory[2087] = 32'h78;
memory[2088] = 32'hf6;
memory[2089] = 32'he7;
memory[2090] = 32'hfe;
memory[2091] = 32'he1;
memory[2092] = 32'hea;
memory[2093] = 32'hfb;
memory[2094] = 32'hf6;
memory[2095] = 32'hf9;
memory[2096] = 32'he6;
memory[2097] = 32'hf9;
memory[2098] = 32'hf6;
memory[2099] = 32'hfb;
memory[2100] = 32'hea;
memory[2101] = 32'he1;
memory[2102] = 32'hfe;
memory[2103] = 32'he7;
memory[2104] = 32'hf6;
memory[2105] = 32'hef;
memory[2106] = 32'hf0;
memory[2107] = 32'hf9;
memory[2108] = 32'hec;
memory[2109] = 32'he7;
memory[2110] = 32'hea;
memory[2111] = 32'hf5;
memory[2112] = 32'hea;
memory[2113] = 32'he7;
memory[2114] = 32'hec;
memory[2115] = 32'hf9;
memory[2116] = 32'hf3;
memory[2117] = 32'hea;
memory[2118] = 32'he9;
memory[2119] = 32'hf0;
memory[2120] = 32'he1;
memory[2121] = 32'hf8;
memory[2122] = 32'hf9;
memory[2123] = 32'he4;
memory[2124] = 32'hf5;
memory[2125] = 32'hf0;
memory[2126] = 32'hf3;
memory[2127] = 32'hfe;
memory[2128] = 32'hf3;
memory[2129] = 32'hf0;
memory[2130] = 32'hf5;
memory[2131] = 32'he4;
memory[2132] = 32'hf9;
memory[2133] = 32'hf8;
memory[2134] = 32'he1;
memory[2135] = 32'hf0;
memory[2136] = 32'he9;
memory[2137] = 32'hea;
memory[2138] = 32'hf3;
memory[2139] = 32'he6;
memory[2140] = 32'he1;
memory[2141] = 32'he4;
memory[2142] = 32'hef;
memory[2143] = 32'he4;
memory[2144] = 32'he1;
memory[2145] = 32'he6;
memory[2146] = 32'h78;
memory[2147] = 32'h78;
memory[2148] = 32'h78;
memory[2149] = 32'h78;
memory[2150] = 32'h78;
memory[2151] = 32'h78;
memory[2152] = 32'hf5;
memory[2153] = 32'he6;
memory[2154] = 32'hfd;
memory[2155] = 32'hfe;
memory[2156] = 32'he9;
memory[2157] = 32'hfa;
memory[2158] = 32'hf5;
memory[2159] = 32'hf8;
memory[2160] = 32'he5;
memory[2161] = 32'hf8;
memory[2162] = 32'hf5;
memory[2163] = 32'hfa;
memory[2164] = 32'he9;
memory[2165] = 32'hfe;
memory[2166] = 32'hfd;
memory[2167] = 32'he6;
memory[2168] = 32'hf5;
memory[2169] = 32'hee;
memory[2170] = 32'hef;
memory[2171] = 32'hf8;
memory[2172] = 32'heb;
memory[2173] = 32'he6;
memory[2174] = 32'he9;
memory[2175] = 32'hf4;
memory[2176] = 32'he9;
memory[2177] = 32'he6;
memory[2178] = 32'heb;
memory[2179] = 32'hf8;
memory[2180] = 32'hf4;
memory[2181] = 32'heb;
memory[2182] = 32'hea;
memory[2183] = 32'hf1;
memory[2184] = 32'he2;
memory[2185] = 32'hf9;
memory[2186] = 32'hfa;
memory[2187] = 32'he5;
memory[2188] = 32'hf6;
memory[2189] = 32'hf1;
memory[2190] = 32'hf4;
memory[2191] = 32'he1;
memory[2192] = 32'hf4;
memory[2193] = 32'hf1;
memory[2194] = 32'hf6;
memory[2195] = 32'he5;
memory[2196] = 32'hfa;
memory[2197] = 32'hf9;
memory[2198] = 32'he2;
memory[2199] = 32'hf1;
memory[2200] = 32'hea;
memory[2201] = 32'heb;
memory[2202] = 32'hf4;
memory[2203] = 32'he7;
memory[2204] = 32'he2;
memory[2205] = 32'he5;
memory[2206] = 32'hf0;
memory[2207] = 32'he5;
memory[2208] = 32'he2;
memory[2209] = 32'he7;
memory[2210] = 32'h78;
memory[2211] = 32'h78;
memory[2212] = 32'h78;
memory[2213] = 32'h78;
memory[2214] = 32'h78;
memory[2215] = 32'h78;
memory[2216] = 32'hf4;
memory[2217] = 32'he5;
memory[2218] = 32'hfc;
memory[2219] = 32'hfd;
memory[2220] = 32'he8;
memory[2221] = 32'hf9;
memory[2222] = 32'hf4;
memory[2223] = 32'hf7;
memory[2224] = 32'he4;
memory[2225] = 32'hf7;
memory[2226] = 32'hf4;
memory[2227] = 32'hf9;
memory[2228] = 32'he8;
memory[2229] = 32'hfd;
memory[2230] = 32'hfc;
memory[2231] = 32'he5;
memory[2232] = 32'hf4;
memory[2233] = 32'hed;
memory[2234] = 32'hee;
memory[2235] = 32'hf7;
memory[2236] = 32'hea;
memory[2237] = 32'he5;
memory[2238] = 32'he8;
memory[2239] = 32'hf3;
memory[2240] = 32'he8;
memory[2241] = 32'he5;
memory[2242] = 32'hea;
memory[2243] = 32'hf7;
memory[2244] = 32'hf5;
memory[2245] = 32'hec;
memory[2246] = 32'heb;
memory[2247] = 32'hf2;
memory[2248] = 32'he3;
memory[2249] = 32'hfa;
memory[2250] = 32'hfb;
memory[2251] = 32'he6;
memory[2252] = 32'hf7;
memory[2253] = 32'hf2;
memory[2254] = 32'hf5;
memory[2255] = 32'he2;
memory[2256] = 32'hf5;
memory[2257] = 32'hf2;
memory[2258] = 32'hf7;
memory[2259] = 32'he6;
memory[2260] = 32'hfb;
memory[2261] = 32'hfa;
memory[2262] = 32'he3;
memory[2263] = 32'hf2;
memory[2264] = 32'heb;
memory[2265] = 32'hec;
memory[2266] = 32'hf5;
memory[2267] = 32'he8;
memory[2268] = 32'he3;
memory[2269] = 32'he6;
memory[2270] = 32'hf1;
memory[2271] = 32'he6;
memory[2272] = 32'he3;
memory[2273] = 32'he5;
memory[2274] = 32'h78;
memory[2275] = 32'h78;
memory[2276] = 32'h78;
memory[2277] = 32'h78;
memory[2278] = 32'h78;
memory[2279] = 32'h78;
memory[2280] = 32'hf3;
memory[2281] = 32'he4;
memory[2282] = 32'hfb;
memory[2283] = 32'hfc;
memory[2284] = 32'he7;
memory[2285] = 32'hf8;
memory[2286] = 32'hf3;
memory[2287] = 32'hf6;
memory[2288] = 32'he3;
memory[2289] = 32'hf6;
memory[2290] = 32'hf3;
memory[2291] = 32'hf8;
memory[2292] = 32'he7;
memory[2293] = 32'hfc;
memory[2294] = 32'hfb;
memory[2295] = 32'he4;
memory[2296] = 32'hf3;
memory[2297] = 32'hec;
memory[2298] = 32'hed;
memory[2299] = 32'hf6;
memory[2300] = 32'he9;
memory[2301] = 32'he4;
memory[2302] = 32'he7;
memory[2303] = 32'hf2;
memory[2304] = 32'he7;
memory[2305] = 32'he4;
memory[2306] = 32'he9;
memory[2307] = 32'hf6;
memory[2308] = 32'hf6;
memory[2309] = 32'hed;
memory[2310] = 32'hec;
memory[2311] = 32'hf3;
memory[2312] = 32'he4;
memory[2313] = 32'hfb;
memory[2314] = 32'hfc;
memory[2315] = 32'he7;
memory[2316] = 32'hf8;
memory[2317] = 32'hf3;
memory[2318] = 32'hf6;
memory[2319] = 32'he3;
memory[2320] = 32'hf6;
memory[2321] = 32'hf3;
memory[2322] = 32'hf8;
memory[2323] = 32'he7;
memory[2324] = 32'hfc;
memory[2325] = 32'hfb;
memory[2326] = 32'he4;
memory[2327] = 32'hf3;
memory[2328] = 32'hec;
memory[2329] = 32'hed;
memory[2330] = 32'hf6;
memory[2331] = 32'he9;
memory[2332] = 32'he4;
memory[2333] = 32'he7;
memory[2334] = 32'hf2;
memory[2335] = 32'he7;
memory[2336] = 32'he9;
memory[2337] = 32'hea;
memory[2338] = 32'h78;
memory[2339] = 32'h78;
memory[2340] = 32'h78;
memory[2341] = 32'h78;
memory[2342] = 32'h78;
memory[2343] = 32'h78;
memory[2344] = 32'hf1;
memory[2345] = 32'he3;
memory[2346] = 32'hfa;
memory[2347] = 32'hfb;
memory[2348] = 32'he6;
memory[2349] = 32'hf7;
memory[2350] = 32'hf2;
memory[2351] = 32'hf5;
memory[2352] = 32'he2;
memory[2353] = 32'hf5;
memory[2354] = 32'hf2;
memory[2355] = 32'hf7;
memory[2356] = 32'he6;
memory[2357] = 32'hfb;
memory[2358] = 32'hfa;
memory[2359] = 32'he3;
memory[2360] = 32'hf2;
memory[2361] = 32'heb;
memory[2362] = 32'hec;
memory[2363] = 32'hf5;
memory[2364] = 32'he8;
memory[2365] = 32'he3;
memory[2366] = 32'he6;
memory[2367] = 32'hf1;
memory[2368] = 32'he6;
memory[2369] = 32'he3;
memory[2370] = 32'he8;
memory[2371] = 32'hf5;
memory[2372] = 32'hf7;
memory[2373] = 32'hee;
memory[2374] = 32'hed;
memory[2375] = 32'hf4;
memory[2376] = 32'he5;
memory[2377] = 32'hfc;
memory[2378] = 32'hfd;
memory[2379] = 32'he8;
memory[2380] = 32'hf9;
memory[2381] = 32'hf4;
memory[2382] = 32'hf7;
memory[2383] = 32'he4;
memory[2384] = 32'hf7;
memory[2385] = 32'hf4;
memory[2386] = 32'hf9;
memory[2387] = 32'he8;
memory[2388] = 32'hfd;
memory[2389] = 32'hfc;
memory[2390] = 32'he5;
memory[2391] = 32'hf4;
memory[2392] = 32'hed;
memory[2393] = 32'hee;
memory[2394] = 32'hf7;
memory[2395] = 32'hea;
memory[2396] = 32'he5;
memory[2397] = 32'he8;
memory[2398] = 32'hf3;
memory[2399] = 32'hf5;
memory[2400] = 32'hf6;
memory[2401] = 32'hf7;
memory[2402] = 32'h78;
memory[2403] = 32'h78;
memory[2404] = 32'h78;
memory[2405] = 32'h65;
memory[2406] = 32'hfc;
memory[2407] = 32'hfd;
memory[2408] = 32'hfe;
memory[2409] = 32'he1;
memory[2410] = 32'hf9;
memory[2411] = 32'hfa;
memory[2412] = 32'he5;
memory[2413] = 32'hf6;
memory[2414] = 32'hf1;
memory[2415] = 32'hf4;
memory[2416] = 32'he1;
memory[2417] = 32'hf4;
memory[2418] = 32'hf1;
memory[2419] = 32'hf6;
memory[2420] = 32'he5;
memory[2421] = 32'hfa;
memory[2422] = 32'hf9;
memory[2423] = 32'he2;
memory[2424] = 32'hf1;
memory[2425] = 32'hea;
memory[2426] = 32'heb;
memory[2427] = 32'hf4;
memory[2428] = 32'he7;
memory[2429] = 32'he2;
memory[2430] = 32'he5;
memory[2431] = 32'hf0;
memory[2432] = 32'he5;
memory[2433] = 32'he2;
memory[2434] = 32'he7;
memory[2435] = 32'hf4;
memory[2436] = 32'hf8;
memory[2437] = 32'hef;
memory[2438] = 32'hee;
memory[2439] = 32'hf5;
memory[2440] = 32'he6;
memory[2441] = 32'hfd;
memory[2442] = 32'hfe;
memory[2443] = 32'he9;
memory[2444] = 32'hfa;
memory[2445] = 32'hf5;
memory[2446] = 32'hf8;
memory[2447] = 32'he5;
memory[2448] = 32'hf8;
memory[2449] = 32'hf5;
memory[2450] = 32'hfa;
memory[2451] = 32'he9;
memory[2452] = 32'hfe;
memory[2453] = 32'hfd;
memory[2454] = 32'he6;
memory[2455] = 32'hf5;
memory[2456] = 32'hee;
memory[2457] = 32'hef;
memory[2458] = 32'hf8;
memory[2459] = 32'heb;
memory[2460] = 32'he6;
memory[2461] = 32'he9;
memory[2462] = 32'heb;
memory[2463] = 32'hec;
memory[2464] = 32'hed;
memory[2465] = 32'hee;
memory[2466] = 32'hef;
memory[2467] = 32'hf0;
memory[2468] = 32'hf1;
memory[2469] = 32'hf2;
memory[2470] = 32'hf3;
memory[2471] = 32'hf4;
memory[2472] = 32'hf5;
memory[2473] = 32'hf6;
memory[2474] = 32'hf7;
memory[2475] = 32'hf9;
memory[2476] = 32'he4;
memory[2477] = 32'hf5;
memory[2478] = 32'hf0;
memory[2479] = 32'hf3;
memory[2480] = 32'hfe;
memory[2481] = 32'hf3;
memory[2482] = 32'hf0;
memory[2483] = 32'hf5;
memory[2484] = 32'he4;
memory[2485] = 32'hf9;
memory[2486] = 32'hf8;
memory[2487] = 32'he1;
memory[2488] = 32'hf0;
memory[2489] = 32'he9;
memory[2490] = 32'hea;
memory[2491] = 32'hf3;
memory[2492] = 32'he6;
memory[2493] = 32'he1;
memory[2494] = 32'he4;
memory[2495] = 32'hef;
memory[2496] = 32'he4;
memory[2497] = 32'he1;
memory[2498] = 32'he6;
memory[2499] = 32'hf3;
memory[2500] = 32'hf9;
memory[2501] = 32'hf0;
memory[2502] = 32'hef;
memory[2503] = 32'hf6;
memory[2504] = 32'he7;
memory[2505] = 32'hfe;
memory[2506] = 32'he1;
memory[2507] = 32'hea;
memory[2508] = 32'hfb;
memory[2509] = 32'hf6;
memory[2510] = 32'hf9;
memory[2511] = 32'he6;
memory[2512] = 32'hf9;
memory[2513] = 32'hf6;
memory[2514] = 32'hfb;
memory[2515] = 32'hea;
memory[2516] = 32'he1;
memory[2517] = 32'hfe;
memory[2518] = 32'he7;
memory[2519] = 32'hf6;
memory[2520] = 32'hef;
memory[2521] = 32'hf0;
memory[2522] = 32'hf9;
memory[2523] = 32'hec;
memory[2524] = 32'he7;
memory[2525] = 32'he9;
memory[2526] = 32'hea;
memory[2527] = 32'heb;
memory[2528] = 32'hec;
memory[2529] = 32'hed;
memory[2530] = 32'hee;
memory[2531] = 32'hef;
memory[2532] = 32'hf0;
memory[2533] = 32'hf1;
memory[2534] = 32'hf2;
memory[2535] = 32'hf3;
memory[2536] = 32'hf4;
memory[2537] = 32'hf5;
memory[2538] = 32'hf6;
memory[2539] = 32'hf7;
memory[2540] = 32'he3;
memory[2541] = 32'hf4;
memory[2542] = 32'hef;
memory[2543] = 32'hf2;
memory[2544] = 32'hfd;
memory[2545] = 32'hf2;
memory[2546] = 32'hef;
memory[2547] = 32'hf4;
memory[2548] = 32'he3;
memory[2549] = 32'hf8;
memory[2550] = 32'hf7;
memory[2551] = 32'hfe;
memory[2552] = 32'hef;
memory[2553] = 32'he8;
memory[2554] = 32'he9;
memory[2555] = 32'hf2;
memory[2556] = 32'he5;
memory[2557] = 32'hfe;
memory[2558] = 32'he3;
memory[2559] = 32'hee;
memory[2560] = 32'he3;
memory[2561] = 32'hfe;
memory[2562] = 32'he5;
memory[2563] = 32'hf2;
memory[2564] = 32'hfa;
memory[2565] = 32'hf1;
memory[2566] = 32'hf0;
memory[2567] = 32'hf7;
memory[2568] = 32'he8;
memory[2569] = 32'he1;
memory[2570] = 32'he2;
memory[2571] = 32'heb;
memory[2572] = 32'hfc;
memory[2573] = 32'hf7;
memory[2574] = 32'hfa;
memory[2575] = 32'he7;
memory[2576] = 32'hfa;
memory[2577] = 32'hf7;
memory[2578] = 32'hfc;
memory[2579] = 32'heb;
memory[2580] = 32'he2;
memory[2581] = 32'he1;
memory[2582] = 32'he8;
memory[2583] = 32'hf7;
memory[2584] = 32'hf0;
memory[2585] = 32'hf1;
memory[2586] = 32'hfa;
memory[2587] = 32'hed;
memory[2588] = 32'hef;
memory[2589] = 32'hf0;
memory[2590] = 32'hf1;
memory[2591] = 32'hf2;
memory[2592] = 32'hf3;
memory[2593] = 32'hf4;
memory[2594] = 32'hf5;
memory[2595] = 32'hf6;
memory[2596] = 32'hf7;
memory[2597] = 32'hf8;
memory[2598] = 32'hf9;
memory[2599] = 32'hfa;
memory[2600] = 32'hfb;
memory[2601] = 32'hfc;
memory[2602] = 32'hfd;
memory[2603] = 32'hfe;
memory[2604] = 32'he1;
memory[2605] = 32'hf3;
memory[2606] = 32'hee;
memory[2607] = 32'hf1;
memory[2608] = 32'hfc;
memory[2609] = 32'hf1;
memory[2610] = 32'hee;
memory[2611] = 32'hf3;
memory[2612] = 32'he2;
memory[2613] = 32'hf7;
memory[2614] = 32'hf6;
memory[2615] = 32'hfd;
memory[2616] = 32'hee;
memory[2617] = 32'he7;
memory[2618] = 32'he8;
memory[2619] = 32'hf1;
memory[2620] = 32'he4;
memory[2621] = 32'hfd;
memory[2622] = 32'he2;
memory[2623] = 32'hed;
memory[2624] = 32'he2;
memory[2625] = 32'hfd;
memory[2626] = 32'he4;
memory[2627] = 32'hf1;
memory[2628] = 32'hfb;
memory[2629] = 32'hf2;
memory[2630] = 32'hf1;
memory[2631] = 32'hf8;
memory[2632] = 32'he9;
memory[2633] = 32'he2;
memory[2634] = 32'he3;
memory[2635] = 32'hec;
memory[2636] = 32'hfd;
memory[2637] = 32'hf8;
memory[2638] = 32'hfb;
memory[2639] = 32'he8;
memory[2640] = 32'hfb;
memory[2641] = 32'hf8;
memory[2642] = 32'hfd;
memory[2643] = 32'hec;
memory[2644] = 32'he3;
memory[2645] = 32'he2;
memory[2646] = 32'he9;
memory[2647] = 32'hf8;
memory[2648] = 32'hf1;
memory[2649] = 32'hf2;
memory[2650] = 32'hfb;
memory[2651] = 32'hfd;
memory[2652] = 32'hfe;
memory[2653] = 32'he1;
memory[2654] = 32'he2;
memory[2655] = 32'he3;
memory[2656] = 32'he4;
memory[2657] = 32'he5;
memory[2658] = 32'he6;
memory[2659] = 32'he7;
memory[2660] = 32'he8;
memory[2661] = 32'he9;
memory[2662] = 32'hea;
memory[2663] = 32'heb;
memory[2664] = 32'hec;
memory[2665] = 32'hed;
memory[2666] = 32'hee;
memory[2667] = 32'hef;
memory[2668] = 32'hf0;
memory[2669] = 32'hf1;
memory[2670] = 32'hed;
memory[2671] = 32'hf0;
memory[2672] = 32'hfb;
memory[2673] = 32'hf0;
memory[2674] = 32'hed;
memory[2675] = 32'hf2;
memory[2676] = 32'he1;
memory[2677] = 32'hf6;
memory[2678] = 32'hf5;
memory[2679] = 32'hfc;
memory[2680] = 32'hed;
memory[2681] = 32'he6;
memory[2682] = 32'he7;
memory[2683] = 32'hf0;
memory[2684] = 32'he3;
memory[2685] = 32'hfc;
memory[2686] = 32'he1;
memory[2687] = 32'hec;
memory[2688] = 32'he1;
memory[2689] = 32'hfc;
memory[2690] = 32'he3;
memory[2691] = 32'hf0;
memory[2692] = 32'hfc;
memory[2693] = 32'hf3;
memory[2694] = 32'hf2;
memory[2695] = 32'hf9;
memory[2696] = 32'hea;
memory[2697] = 32'he3;
memory[2698] = 32'he4;
memory[2699] = 32'hed;
memory[2700] = 32'hfe;
memory[2701] = 32'hf9;
memory[2702] = 32'hfc;
memory[2703] = 32'he9;
memory[2704] = 32'hfc;
memory[2705] = 32'hf9;
memory[2706] = 32'hfe;
memory[2707] = 32'hed;
memory[2708] = 32'he4;
memory[2709] = 32'he3;
memory[2710] = 32'hea;
memory[2711] = 32'hf9;
memory[2712] = 32'hf2;
memory[2713] = 32'hf3;
memory[2714] = 32'hf5;
memory[2715] = 32'hf6;
memory[2716] = 32'hf7;
memory[2717] = 32'hf8;
memory[2718] = 32'hf9;
memory[2719] = 32'hfa;
memory[2720] = 32'hfb;
memory[2721] = 32'hfc;
memory[2722] = 32'hfd;
memory[2723] = 32'hfe;
memory[2724] = 32'he1;
memory[2725] = 32'he2;
memory[2726] = 32'he3;
memory[2727] = 32'he4;
memory[2728] = 32'he5;
memory[2729] = 32'he6;
memory[2730] = 32'he7;
memory[2731] = 32'he8;
memory[2732] = 32'he9;
memory[2733] = 32'hea;
memory[2734] = 32'heb;
memory[2735] = 32'hef;
memory[2736] = 32'hfa;
memory[2737] = 32'hef;
memory[2738] = 32'hec;
memory[2739] = 32'hf1;
memory[2740] = 32'hfe;
memory[2741] = 32'hf5;
memory[2742] = 32'hf4;
memory[2743] = 32'hfb;
memory[2744] = 32'hec;
memory[2745] = 32'he5;
memory[2746] = 32'he6;
memory[2747] = 32'hef;
memory[2748] = 32'he2;
memory[2749] = 32'hfb;
memory[2750] = 32'hfe;
memory[2751] = 32'heb;
memory[2752] = 32'hfe;
memory[2753] = 32'hfb;
memory[2754] = 32'he2;
memory[2755] = 32'hef;
memory[2756] = 32'hfd;
memory[2757] = 32'hf4;
memory[2758] = 32'hf3;
memory[2759] = 32'hfa;
memory[2760] = 32'heb;
memory[2761] = 32'he4;
memory[2762] = 32'he5;
memory[2763] = 32'hee;
memory[2764] = 32'he1;
memory[2765] = 32'hfa;
memory[2766] = 32'hfd;
memory[2767] = 32'hea;
memory[2768] = 32'hfd;
memory[2769] = 32'hfa;
memory[2770] = 32'he1;
memory[2771] = 32'hee;
memory[2772] = 32'he5;
memory[2773] = 32'he4;
memory[2774] = 32'heb;
memory[2775] = 32'hfa;
memory[2776] = 32'hf3;
memory[2777] = 32'hf5;
memory[2778] = 32'hf6;
memory[2779] = 32'hf7;
memory[2780] = 32'hf8;
memory[2781] = 32'hf9;
memory[2782] = 32'hfa;
memory[2783] = 32'hfb;
memory[2784] = 32'hfc;
memory[2785] = 32'hfd;
memory[2786] = 32'hfe;
memory[2787] = 32'he1;
memory[2788] = 32'he2;
memory[2789] = 32'he3;
memory[2790] = 32'he4;
memory[2791] = 32'he5;
memory[2792] = 32'he6;
memory[2793] = 32'he7;
memory[2794] = 32'he8;
memory[2795] = 32'he9;
memory[2796] = 32'hea;
memory[2797] = 32'heb;
memory[2798] = 32'hec;
memory[2799] = 32'hed;
memory[2800] = 32'hf9;
memory[2801] = 32'hee;
memory[2802] = 32'heb;
memory[2803] = 32'hf0;
memory[2804] = 32'hfd;
memory[2805] = 32'hf4;
memory[2806] = 32'hf3;
memory[2807] = 32'hfa;
memory[2808] = 32'heb;
memory[2809] = 32'he4;
memory[2810] = 32'he5;
memory[2811] = 32'hee;
memory[2812] = 32'he1;
memory[2813] = 32'hfa;
memory[2814] = 32'hfd;
memory[2815] = 32'hea;
memory[2816] = 32'hfd;
memory[2817] = 32'hfa;
memory[2818] = 32'he1;
memory[2819] = 32'hee;
memory[2820] = 32'hfe;
memory[2821] = 32'hf5;
memory[2822] = 32'hf4;
memory[2823] = 32'hfb;
memory[2824] = 32'hec;
memory[2825] = 32'he5;
memory[2826] = 32'he6;
memory[2827] = 32'hef;
memory[2828] = 32'he2;
memory[2829] = 32'hfb;
memory[2830] = 32'hfe;
memory[2831] = 32'heb;
memory[2832] = 32'hfe;
memory[2833] = 32'hfb;
memory[2834] = 32'he2;
memory[2835] = 32'hef;
memory[2836] = 32'he6;
memory[2837] = 32'he5;
memory[2838] = 32'hec;
memory[2839] = 32'hfb;
memory[2840] = 32'hfd;
memory[2841] = 32'hfe;
memory[2842] = 32'he1;
memory[2843] = 32'he2;
memory[2844] = 32'he3;
memory[2845] = 32'he4;
memory[2846] = 32'he5;
memory[2847] = 32'he6;
memory[2848] = 32'he7;
memory[2849] = 32'he8;
memory[2850] = 32'he9;
memory[2851] = 32'hea;
memory[2852] = 32'heb;
memory[2853] = 32'hec;
memory[2854] = 32'hed;
memory[2855] = 32'hee;
memory[2856] = 32'hef;
memory[2857] = 32'hf0;
memory[2858] = 32'hf1;
memory[2859] = 32'hf2;
memory[2860] = 32'hf3;
memory[2861] = 32'hf4;
memory[2862] = 32'hf5;
memory[2863] = 32'hf6;
memory[2864] = 32'hf7;
memory[2865] = 32'hed;
memory[2866] = 32'hea;
memory[2867] = 32'hef;
memory[2868] = 32'hfc;
memory[2869] = 32'hf3;
memory[2870] = 32'hf2;
memory[2871] = 32'hf9;
memory[2872] = 32'hea;
memory[2873] = 32'he3;
memory[2874] = 32'he4;
memory[2875] = 32'hed;
memory[2876] = 32'hfe;
memory[2877] = 32'hf9;
memory[2878] = 32'hfc;
memory[2879] = 32'he9;
memory[2880] = 32'hfc;
memory[2881] = 32'hf9;
memory[2882] = 32'hfe;
memory[2883] = 32'hed;
memory[2884] = 32'he1;
memory[2885] = 32'hf6;
memory[2886] = 32'hf5;
memory[2887] = 32'hfc;
memory[2888] = 32'hed;
memory[2889] = 32'he6;
memory[2890] = 32'he7;
memory[2891] = 32'hf0;
memory[2892] = 32'he3;
memory[2893] = 32'hfc;
memory[2894] = 32'he1;
memory[2895] = 32'hec;
memory[2896] = 32'he1;
memory[2897] = 32'hfc;
memory[2898] = 32'he3;
memory[2899] = 32'hf0;
memory[2900] = 32'he7;
memory[2901] = 32'he6;
memory[2902] = 32'hed;
memory[2903] = 32'hef;
memory[2904] = 32'hf0;
memory[2905] = 32'hf1;
memory[2906] = 32'hf2;
memory[2907] = 32'hf3;
memory[2908] = 32'hf4;
memory[2909] = 32'hf5;
memory[2910] = 32'hf6;
memory[2911] = 32'hf7;
memory[2912] = 32'hf8;
memory[2913] = 32'hf9;
memory[2914] = 32'hfa;
memory[2915] = 32'hfb;
memory[2916] = 32'hfc;
memory[2917] = 32'hfd;
memory[2918] = 32'hfe;
memory[2919] = 32'he1;
memory[2920] = 32'he2;
memory[2921] = 32'he3;
memory[2922] = 32'he4;
memory[2923] = 32'he5;
memory[2924] = 32'he6;
memory[2925] = 32'he7;
memory[2926] = 32'he8;
memory[2927] = 32'he9;
memory[2928] = 32'hea;
memory[2929] = 32'heb;
memory[2930] = 32'he9;
memory[2931] = 32'hee;
memory[2932] = 32'hfb;
memory[2933] = 32'hf2;
memory[2934] = 32'hf1;
memory[2935] = 32'hf8;
memory[2936] = 32'he9;
memory[2937] = 32'he2;
memory[2938] = 32'he3;
memory[2939] = 32'hec;
memory[2940] = 32'hfd;
memory[2941] = 32'hf8;
memory[2942] = 32'hfb;
memory[2943] = 32'he8;
memory[2944] = 32'hfb;
memory[2945] = 32'hf8;
memory[2946] = 32'hfd;
memory[2947] = 32'hec;
memory[2948] = 32'he2;
memory[2949] = 32'hf7;
memory[2950] = 32'hf6;
memory[2951] = 32'hfd;
memory[2952] = 32'hee;
memory[2953] = 32'he7;
memory[2954] = 32'he8;
memory[2955] = 32'hf1;
memory[2956] = 32'he4;
memory[2957] = 32'hfd;
memory[2958] = 32'he2;
memory[2959] = 32'hed;
memory[2960] = 32'he2;
memory[2961] = 32'hfd;
memory[2962] = 32'he4;
memory[2963] = 32'hf1;
memory[2964] = 32'he8;
memory[2965] = 32'he7;
memory[2966] = 32'he9;
memory[2967] = 32'hea;
memory[2968] = 32'heb;
memory[2969] = 32'hec;
memory[2970] = 32'hed;
memory[2971] = 32'hee;
memory[2972] = 32'hef;
memory[2973] = 32'hf0;
memory[2974] = 32'hf1;
memory[2975] = 32'hf2;
memory[2976] = 32'hf3;
memory[2977] = 32'hf4;
memory[2978] = 32'hf5;
memory[2979] = 32'hf6;
memory[2980] = 32'hf7;
memory[2981] = 32'hf8;
memory[2982] = 32'hf9;
memory[2983] = 32'hfa;
memory[2984] = 32'hfb;
memory[2985] = 32'hfc;
memory[2986] = 32'hfd;
memory[2987] = 32'hfe;
memory[2988] = 32'he1;
memory[2989] = 32'he2;
memory[2990] = 32'he3;
memory[2991] = 32'he4;
memory[2992] = 32'he5;
memory[2993] = 32'he6;
memory[2994] = 32'he7;
memory[2995] = 32'hed;
memory[2996] = 32'hfa;
memory[2997] = 32'hf1;
memory[2998] = 32'hf0;
memory[2999] = 32'hf7;
memory[3000] = 32'he8;
memory[3001] = 32'he1;
memory[3002] = 32'he2;
memory[3003] = 32'heb;
memory[3004] = 32'hfc;
memory[3005] = 32'hf7;
memory[3006] = 32'hfa;
memory[3007] = 32'he7;
memory[3008] = 32'hfa;
memory[3009] = 32'hf7;
memory[3010] = 32'hfc;
memory[3011] = 32'heb;
memory[3012] = 32'he3;
memory[3013] = 32'hf8;
memory[3014] = 32'hf7;
memory[3015] = 32'hfe;
memory[3016] = 32'hef;
memory[3017] = 32'he8;
memory[3018] = 32'he9;
memory[3019] = 32'hf2;
memory[3020] = 32'he5;
memory[3021] = 32'hfe;
memory[3022] = 32'he3;
memory[3023] = 32'hee;
memory[3024] = 32'he3;
memory[3025] = 32'hfe;
memory[3026] = 32'he5;
memory[3027] = 32'hf2;
memory[3028] = 32'he9;
memory[3029] = 32'heb;
memory[3030] = 32'hec;
memory[3031] = 32'hed;
memory[3032] = 32'hee;
memory[3033] = 32'hef;
memory[3034] = 32'hf0;
memory[3035] = 32'hf1;
memory[3036] = 32'hf2;
memory[3037] = 32'hf3;
memory[3038] = 32'hf4;
memory[3039] = 32'hf5;
memory[3040] = 32'hf6;
memory[3041] = 32'hf7;
memory[3042] = 32'hf8;
memory[3043] = 32'hf9;
memory[3044] = 32'hfa;
memory[3045] = 32'hfb;
memory[3046] = 32'hfc;
memory[3047] = 32'hfd;
memory[3048] = 32'hfe;
memory[3049] = 32'he1;
memory[3050] = 32'he2;
memory[3051] = 32'he3;
memory[3052] = 32'he4;
memory[3053] = 32'he5;
memory[3054] = 32'he6;
memory[3055] = 32'he7;
memory[3056] = 32'he8;
memory[3057] = 32'he9;
memory[3058] = 32'hea;
memory[3059] = 32'heb;
memory[3060] = 32'hf9;
memory[3061] = 32'hf0;
memory[3062] = 32'hef;
memory[3063] = 32'hf6;
memory[3064] = 32'he7;
memory[3065] = 32'hfe;
memory[3066] = 32'he1;
memory[3067] = 32'hea;
memory[3068] = 32'hfb;
memory[3069] = 32'hf6;
memory[3070] = 32'hf9;
memory[3071] = 32'he6;
memory[3072] = 32'hf9;
memory[3073] = 32'hf6;
memory[3074] = 32'hfb;
memory[3075] = 32'hea;
memory[3076] = 32'he4;
memory[3077] = 32'hf9;
memory[3078] = 32'hf8;
memory[3079] = 32'he1;
memory[3080] = 32'hf0;
memory[3081] = 32'he9;
memory[3082] = 32'hea;
memory[3083] = 32'hf3;
memory[3084] = 32'he6;
memory[3085] = 32'he1;
memory[3086] = 32'he4;
memory[3087] = 32'hef;
memory[3088] = 32'he4;
memory[3089] = 32'he1;
memory[3090] = 32'he6;
memory[3091] = 32'hf3;
memory[3092] = 32'hf5;
memory[3093] = 32'hf6;
memory[3094] = 32'hf7;
memory[3095] = 32'hf8;
memory[3096] = 32'hf9;
memory[3097] = 32'hfa;
memory[3098] = 32'hfb;
memory[3099] = 32'hfc;
memory[3100] = 32'hfd;
memory[3101] = 32'hfe;
memory[3102] = 32'he1;
memory[3103] = 32'he2;
memory[3104] = 32'he3;
memory[3105] = 32'he4;
memory[3106] = 32'he5;
memory[3107] = 32'he6;
memory[3108] = 32'he7;
memory[3109] = 32'he8;
memory[3110] = 32'he9;
memory[3111] = 32'hea;
memory[3112] = 32'heb;
memory[3113] = 32'hec;
memory[3114] = 32'hed;
memory[3115] = 32'hee;
memory[3116] = 32'hef;
memory[3117] = 32'hf0;
memory[3118] = 32'hf1;
memory[3119] = 32'hf2;
memory[3120] = 32'hf3;
memory[3121] = 32'hf4;
memory[3122] = 32'hf5;
memory[3123] = 32'hf6;
memory[3124] = 32'hf7;
memory[3125] = 32'hef;
memory[3126] = 32'hee;
memory[3127] = 32'hf5;
memory[3128] = 32'he6;
memory[3129] = 32'hfd;
memory[3130] = 32'hfe;
memory[3131] = 32'he9;
memory[3132] = 32'hfa;
memory[3133] = 32'hf5;
memory[3134] = 32'hf8;
memory[3135] = 32'he5;
memory[3136] = 32'hf8;
memory[3137] = 32'hf5;
memory[3138] = 32'hfa;
memory[3139] = 32'he9;
memory[3140] = 32'he5;
memory[3141] = 32'hfa;
memory[3142] = 32'hf9;
memory[3143] = 32'he2;
memory[3144] = 32'hf1;
memory[3145] = 32'hea;
memory[3146] = 32'heb;
memory[3147] = 32'hf4;
memory[3148] = 32'he7;
memory[3149] = 32'he2;
memory[3150] = 32'he5;
memory[3151] = 32'hf0;
memory[3152] = 32'he5;
memory[3153] = 32'he2;
memory[3154] = 32'he7;
memory[3155] = 32'he9;
memory[3156] = 32'hea;
memory[3157] = 32'heb;
memory[3158] = 32'hec;
memory[3159] = 32'hed;
memory[3160] = 32'hee;
memory[3161] = 32'hef;
memory[3162] = 32'hf0;
memory[3163] = 32'hf1;
memory[3164] = 32'hf2;
memory[3165] = 32'hf3;
memory[3166] = 32'hf4;
memory[3167] = 32'hf5;
memory[3168] = 32'hf6;
memory[3169] = 32'hf7;
memory[3170] = 32'hf8;
memory[3171] = 32'hf9;
memory[3172] = 32'hfa;
memory[3173] = 32'hfb;
memory[3174] = 32'hfc;
memory[3175] = 32'hfd;
memory[3176] = 32'hfe;
memory[3177] = 32'he1;
memory[3178] = 32'he2;
memory[3179] = 32'he3;
memory[3180] = 32'he4;
memory[3181] = 32'he5;
memory[3182] = 32'he6;
memory[3183] = 32'he7;
memory[3184] = 32'he8;
memory[3185] = 32'he9;
memory[3186] = 32'hea;
memory[3187] = 32'heb;
memory[3188] = 32'hec;
memory[3189] = 32'hed;
memory[3190] = 32'hed;
memory[3191] = 32'hf4;
memory[3192] = 32'he5;
memory[3193] = 32'hfc;
memory[3194] = 32'hfd;
memory[3195] = 32'he8;
memory[3196] = 32'hf9;
memory[3197] = 32'hf4;
memory[3198] = 32'hf7;
memory[3199] = 32'he4;
memory[3200] = 32'hf7;
memory[3201] = 32'hf4;
memory[3202] = 32'hf9;
memory[3203] = 32'he8;
memory[3204] = 32'he6;
memory[3205] = 32'hfb;
memory[3206] = 32'hfa;
memory[3207] = 32'he3;
memory[3208] = 32'hf2;
memory[3209] = 32'heb;
memory[3210] = 32'hec;
memory[3211] = 32'hf5;
memory[3212] = 32'he8;
memory[3213] = 32'he3;
memory[3214] = 32'he6;
memory[3215] = 32'hf1;
memory[3216] = 32'he6;
memory[3217] = 32'he3;
memory[3218] = 32'he5;
memory[3219] = 32'he6;
memory[3220] = 32'he7;
memory[3221] = 32'he8;
memory[3222] = 32'he9;
memory[3223] = 32'hea;
memory[3224] = 32'heb;
memory[3225] = 32'hec;
memory[3226] = 32'hed;
memory[3227] = 32'hee;
memory[3228] = 32'hef;
memory[3229] = 32'hf0;
memory[3230] = 32'hf1;
memory[3231] = 32'hf2;
memory[3232] = 32'hf3;
memory[3233] = 32'hf4;
memory[3234] = 32'hf5;
memory[3235] = 32'hf6;
memory[3236] = 32'hf7;
memory[3237] = 32'hf8;
memory[3238] = 32'hf9;
memory[3239] = 32'hfa;
memory[3240] = 32'hfb;
memory[3241] = 32'hfc;
memory[3242] = 32'hfd;
memory[3243] = 32'hfe;
memory[3244] = 32'he1;
memory[3245] = 32'he2;
memory[3246] = 32'he3;
memory[3247] = 32'he4;
memory[3248] = 32'he5;
memory[3249] = 32'he6;
memory[3250] = 32'he7;
memory[3251] = 32'he8;
memory[3252] = 32'he9;
memory[3253] = 32'hea;
memory[3254] = 32'heb;
memory[3255] = 32'hf3;
memory[3256] = 32'h66;
memory[3257] = 32'h66;
memory[3258] = 32'h66;
memory[3259] = 32'h66;
memory[3260] = 32'hf8;
memory[3261] = 32'hf3;
memory[3262] = 32'hf6;
memory[3263] = 32'he3;
memory[3264] = 32'hf6;
memory[3265] = 32'hf3;
memory[3266] = 32'hf8;
memory[3267] = 32'he7;
memory[3268] = 32'he7;
memory[3269] = 32'hfc;
memory[3270] = 32'hfb;
memory[3271] = 32'he4;
memory[3272] = 32'hf3;
memory[3273] = 32'hec;
memory[3274] = 32'hed;
memory[3275] = 32'hf6;
memory[3276] = 32'he9;
memory[3277] = 32'he4;
memory[3278] = 32'he7;
memory[3279] = 32'hf2;
memory[3280] = 32'he7;
memory[3281] = 32'he9;
memory[3282] = 32'hea;
memory[3283] = 32'heb;
memory[3284] = 32'hec;
memory[3285] = 32'hed;
memory[3286] = 32'hee;
memory[3287] = 32'hef;
memory[3288] = 32'hf0;
memory[3289] = 32'hf1;
memory[3290] = 32'hf2;
memory[3291] = 32'hf3;
memory[3292] = 32'hf4;
memory[3293] = 32'hf5;
memory[3294] = 32'hf6;
memory[3295] = 32'hf7;
memory[3296] = 32'hf8;
memory[3297] = 32'hf9;
memory[3298] = 32'hfa;
memory[3299] = 32'hfb;
memory[3300] = 32'hfc;
memory[3301] = 32'hfd;
memory[3302] = 32'hfe;
memory[3303] = 32'he1;
memory[3304] = 32'he2;
memory[3305] = 32'he3;
memory[3306] = 32'he4;
memory[3307] = 32'he5;
memory[3308] = 32'he6;
memory[3309] = 32'he7;
memory[3310] = 32'he8;
memory[3311] = 32'he9;
memory[3312] = 32'hea;
memory[3313] = 32'heb;
memory[3314] = 32'hec;
memory[3315] = 32'hed;
memory[3316] = 32'hee;
memory[3317] = 32'hef;
memory[3318] = 32'hf0;
memory[3319] = 32'hf1;
memory[3320] = 32'h66;
memory[3321] = 32'h66;
memory[3322] = 32'h66;
memory[3323] = 32'h66;
memory[3324] = 32'hf7;
memory[3325] = 32'hf2;
memory[3326] = 32'hf5;
memory[3327] = 32'he2;
memory[3328] = 32'hf5;
memory[3329] = 32'hf2;
memory[3330] = 32'hf7;
memory[3331] = 32'he6;
memory[3332] = 32'he8;
memory[3333] = 32'hfd;
memory[3334] = 32'hfc;
memory[3335] = 32'he5;
memory[3336] = 32'hf4;
memory[3337] = 32'hed;
memory[3338] = 32'hee;
memory[3339] = 32'hf7;
memory[3340] = 32'hea;
memory[3341] = 32'he5;
memory[3342] = 32'he8;
memory[3343] = 32'hf3;
memory[3344] = 32'hf5;
memory[3345] = 32'hf6;
memory[3346] = 32'hf7;
memory[3347] = 32'hf8;
memory[3348] = 32'hf9;
memory[3349] = 32'hfa;
memory[3350] = 32'hfb;
memory[3351] = 32'hfc;
memory[3352] = 32'hfd;
memory[3353] = 32'hfe;
memory[3354] = 32'he1;
memory[3355] = 32'he2;
memory[3356] = 32'he3;
memory[3357] = 32'he4;
memory[3358] = 32'he5;
memory[3359] = 32'he6;
memory[3360] = 32'he7;
memory[3361] = 32'he8;
memory[3362] = 32'he9;
memory[3363] = 32'hea;
memory[3364] = 32'heb;
memory[3365] = 32'hec;
memory[3366] = 32'hed;
memory[3367] = 32'hee;
memory[3368] = 32'hef;
memory[3369] = 32'hf0;
memory[3370] = 32'hf1;
memory[3371] = 32'hf2;
memory[3372] = 32'hf3;
memory[3373] = 32'hf4;
memory[3374] = 32'hf5;
memory[3375] = 32'hf6;
memory[3376] = 32'hf7;
memory[3377] = 32'hf8;
memory[3378] = 32'hf9;
memory[3379] = 32'hfa;
memory[3380] = 32'hfb;
memory[3381] = 32'hfc;
memory[3382] = 32'hfd;
memory[3383] = 32'hfe;
memory[3384] = 32'h66;
memory[3385] = 32'h66;
memory[3386] = 32'h66;
memory[3387] = 32'h66;
memory[3388] = 32'hf6;
memory[3389] = 32'hf1;
memory[3390] = 32'hf4;
memory[3391] = 32'he1;
memory[3392] = 32'hf4;
memory[3393] = 32'hf1;
memory[3394] = 32'hf6;
memory[3395] = 32'he5;
memory[3396] = 32'he9;
memory[3397] = 32'hfe;
memory[3398] = 32'hfd;
memory[3399] = 32'he6;
memory[3400] = 32'hf5;
memory[3401] = 32'hee;
memory[3402] = 32'hef;
memory[3403] = 32'hf8;
memory[3404] = 32'heb;
memory[3405] = 32'he6;
memory[3406] = 32'he9;
memory[3407] = 32'heb;
memory[3408] = 32'hec;
memory[3409] = 32'hed;
memory[3410] = 32'hee;
memory[3411] = 32'hef;
memory[3412] = 32'hf0;
memory[3413] = 32'hf1;
memory[3414] = 32'hf2;
memory[3415] = 32'hf3;
memory[3416] = 32'hf4;
memory[3417] = 32'hf5;
memory[3418] = 32'hf6;
memory[3419] = 32'hf7;
memory[3420] = 32'hf8;
memory[3421] = 32'hf9;
memory[3422] = 32'hfa;
memory[3423] = 32'hfb;
memory[3424] = 32'hfc;
memory[3425] = 32'hfd;
memory[3426] = 32'hfe;
memory[3427] = 32'he1;
memory[3428] = 32'he2;
memory[3429] = 32'he3;
memory[3430] = 32'he4;
memory[3431] = 32'he5;
memory[3432] = 32'he6;
memory[3433] = 32'he7;
memory[3434] = 32'he8;
memory[3435] = 32'he9;
memory[3436] = 32'hea;
memory[3437] = 32'heb;
memory[3438] = 32'hec;
memory[3439] = 32'hed;
memory[3440] = 32'hee;
memory[3441] = 32'hef;
memory[3442] = 32'hf0;
memory[3443] = 32'hf1;
memory[3444] = 32'hf2;
memory[3445] = 32'hf3;
memory[3446] = 32'hf4;
memory[3447] = 32'hf5;
memory[3448] = 32'h66;
memory[3449] = 32'h66;
memory[3450] = 32'h66;
memory[3451] = 32'h66;
memory[3452] = 32'hf5;
memory[3453] = 32'hf0;
memory[3454] = 32'hf3;
memory[3455] = 32'hfe;
memory[3456] = 32'hf3;
memory[3457] = 32'hf0;
memory[3458] = 32'hf5;
memory[3459] = 32'he4;
memory[3460] = 32'hea;
memory[3461] = 32'he1;
memory[3462] = 32'hfe;
memory[3463] = 32'he7;
memory[3464] = 32'hf6;
memory[3465] = 32'hef;
memory[3466] = 32'hf0;
memory[3467] = 32'hf9;
memory[3468] = 32'hec;
memory[3469] = 32'he7;
memory[3470] = 32'he9;
memory[3471] = 32'hea;
memory[3472] = 32'heb;
memory[3473] = 32'hec;
memory[3474] = 32'hed;
memory[3475] = 32'hee;
memory[3476] = 32'hef;
memory[3477] = 32'hf0;
memory[3478] = 32'hf1;
memory[3479] = 32'hf2;
memory[3480] = 32'hf3;
memory[3481] = 32'hf4;
memory[3482] = 32'hf5;
memory[3483] = 32'hf6;
memory[3484] = 32'hf7;
memory[3485] = 32'hf8;
memory[3486] = 32'hf9;
memory[3487] = 32'hfa;
memory[3488] = 32'hfb;
memory[3489] = 32'hfc;
memory[3490] = 32'hfd;
memory[3491] = 32'hfe;
memory[3492] = 32'he1;
memory[3493] = 32'he2;
memory[3494] = 32'he3;
memory[3495] = 32'he4;
memory[3496] = 32'he5;
memory[3497] = 32'he6;
memory[3498] = 32'he7;
memory[3499] = 32'he8;
memory[3500] = 32'he9;
memory[3501] = 32'hea;
memory[3502] = 32'heb;
memory[3503] = 32'hec;
memory[3504] = 32'hed;
memory[3505] = 32'hee;
memory[3506] = 32'hef;
memory[3507] = 32'hf0;
memory[3508] = 32'hf1;
memory[3509] = 32'hf2;
memory[3510] = 32'hf3;
memory[3511] = 32'hf4;
memory[3512] = 32'hf5;
memory[3513] = 32'hf6;
memory[3514] = 32'hf7;
memory[3515] = 32'he3;
memory[3516] = 32'hf4;
memory[3517] = 32'hef;
memory[3518] = 32'hf2;
memory[3519] = 32'hfd;
memory[3520] = 32'hf2;
memory[3521] = 32'hef;
memory[3522] = 32'hf4;
memory[3523] = 32'he3;
memory[3524] = 32'heb;
memory[3525] = 32'he2;
memory[3526] = 32'he1;
memory[3527] = 32'he8;
memory[3528] = 32'hf7;
memory[3529] = 32'hf0;
memory[3530] = 32'hf1;
memory[3531] = 32'hfa;
memory[3532] = 32'hed;
memory[3533] = 32'hef;
memory[3534] = 32'hf0;
memory[3535] = 32'hf1;
memory[3536] = 32'hf2;
memory[3537] = 32'hf3;
memory[3538] = 32'hf4;
memory[3539] = 32'hf5;
memory[3540] = 32'hf6;
memory[3541] = 32'hf7;
memory[3542] = 32'hf8;
memory[3543] = 32'hf9;
memory[3544] = 32'hfa;
memory[3545] = 32'hfb;
memory[3546] = 32'hfc;
memory[3547] = 32'hfd;
memory[3548] = 32'hfe;
memory[3549] = 32'he1;
memory[3550] = 32'he2;
memory[3551] = 32'he3;
memory[3552] = 32'he4;
memory[3553] = 32'he5;
memory[3554] = 32'he6;
memory[3555] = 32'he7;
memory[3556] = 32'he8;
memory[3557] = 32'he9;
memory[3558] = 32'hea;
memory[3559] = 32'heb;
memory[3560] = 32'hec;
memory[3561] = 32'hed;
memory[3562] = 32'hee;
memory[3563] = 32'hef;
memory[3564] = 32'hf0;
memory[3565] = 32'hf1;
memory[3566] = 32'hf2;
memory[3567] = 32'hf3;
memory[3568] = 32'hf4;
memory[3569] = 32'hf5;
memory[3570] = 32'hf6;
memory[3571] = 32'hf7;
memory[3572] = 32'hf8;
memory[3573] = 32'hf9;
memory[3574] = 32'hfa;
memory[3575] = 32'hfb;
memory[3576] = 32'hfc;
memory[3577] = 32'hfd;
memory[3578] = 32'hfe;
memory[3579] = 32'he1;
memory[3580] = 32'hf3;
memory[3581] = 32'hee;
memory[3582] = 32'hf1;
memory[3583] = 32'hfc;
memory[3584] = 32'hf1;
memory[3585] = 32'hee;
memory[3586] = 32'hf3;
memory[3587] = 32'he2;
memory[3588] = 32'hec;
memory[3589] = 32'he3;
memory[3590] = 32'he2;
memory[3591] = 32'he9;
memory[3592] = 32'hf8;
memory[3593] = 32'hf1;
memory[3594] = 32'hf2;
memory[3595] = 32'hfb;
memory[3596] = 32'hfd;
memory[3597] = 32'hfe;
memory[3598] = 32'he1;
memory[3599] = 32'he2;
memory[3600] = 32'he3;
memory[3601] = 32'he4;
memory[3602] = 32'he5;
memory[3603] = 32'he6;
memory[3604] = 32'he7;
memory[3605] = 32'he8;
memory[3606] = 32'he9;
memory[3607] = 32'hea;
memory[3608] = 32'heb;
memory[3609] = 32'hec;
memory[3610] = 32'hed;
memory[3611] = 32'hee;
memory[3612] = 32'hef;
memory[3613] = 32'hf0;
memory[3614] = 32'hf1;
memory[3615] = 32'hf2;
memory[3616] = 32'hf3;
memory[3617] = 32'hf4;
memory[3618] = 32'hf5;
memory[3619] = 32'hf6;
memory[3620] = 32'hf7;
memory[3621] = 32'hf8;
memory[3622] = 32'hf9;
memory[3623] = 32'hfa;
memory[3624] = 32'hfb;
memory[3625] = 32'hfc;
memory[3626] = 32'hfd;
memory[3627] = 32'hfe;
memory[3628] = 32'he1;
memory[3629] = 32'he2;
memory[3630] = 32'he3;
memory[3631] = 32'he4;
memory[3632] = 32'he5;
memory[3633] = 32'he6;
memory[3634] = 32'he7;
memory[3635] = 32'he8;
memory[3636] = 32'he9;
memory[3637] = 32'hea;
memory[3638] = 32'heb;
memory[3639] = 32'hec;
memory[3640] = 32'hed;
memory[3641] = 32'hee;
memory[3642] = 32'hef;
memory[3643] = 32'hf0;
memory[3644] = 32'hf1;
memory[3645] = 32'hed;
memory[3646] = 32'hf0;
memory[3647] = 32'hfb;
memory[3648] = 32'hf0;
memory[3649] = 32'hed;
memory[3650] = 32'hf2;
memory[3651] = 32'he1;
memory[3652] = 32'hed;
memory[3653] = 32'he4;
memory[3654] = 32'he3;
memory[3655] = 32'hea;
memory[3656] = 32'hf9;
memory[3657] = 32'hf2;
memory[3658] = 32'hf3;
memory[3659] = 32'hf5;
memory[3660] = 32'hf6;
memory[3661] = 32'hf7;
memory[3662] = 32'hf8;
memory[3663] = 32'hf9;
memory[3664] = 32'hfa;
memory[3665] = 32'hfb;
memory[3666] = 32'hfc;
memory[3667] = 32'hfd;
memory[3668] = 32'hfe;
memory[3669] = 32'he1;
memory[3670] = 32'he2;
memory[3671] = 32'he3;
memory[3672] = 32'he4;
memory[3673] = 32'he5;
memory[3674] = 32'he6;
memory[3675] = 32'he7;
memory[3676] = 32'he8;
memory[3677] = 32'he9;
memory[3678] = 32'hea;
memory[3679] = 32'heb;
memory[3680] = 32'hec;
memory[3681] = 32'hed;
memory[3682] = 32'hee;
memory[3683] = 32'hef;
memory[3684] = 32'hf0;
memory[3685] = 32'hf1;
memory[3686] = 32'hf2;
memory[3687] = 32'hf3;
memory[3688] = 32'hf4;
memory[3689] = 32'hf5;
memory[3690] = 32'hf6;
memory[3691] = 32'hf7;
memory[3692] = 32'hf8;
memory[3693] = 32'hf9;
memory[3694] = 32'hfa;
memory[3695] = 32'hfb;
memory[3696] = 32'hfc;
memory[3697] = 32'hfd;
memory[3698] = 32'hfe;
memory[3699] = 32'he1;
memory[3700] = 32'he2;
memory[3701] = 32'he3;
memory[3702] = 32'he4;
memory[3703] = 32'he5;
memory[3704] = 32'he6;
memory[3705] = 32'he7;
memory[3706] = 32'he8;
memory[3707] = 32'he9;
memory[3708] = 32'hea;
memory[3709] = 32'heb;
memory[3710] = 32'hef;
memory[3711] = 32'hfa;
memory[3712] = 32'hef;
memory[3713] = 32'hec;
memory[3714] = 32'hf1;
memory[3715] = 32'hfe;
memory[3716] = 32'hee;
memory[3717] = 32'he5;
memory[3718] = 32'he4;
memory[3719] = 32'heb;
memory[3720] = 32'hfa;
memory[3721] = 32'hf3;
memory[3722] = 32'hf5;
memory[3723] = 32'hf6;
memory[3724] = 32'hf7;
memory[3725] = 32'hf8;
memory[3726] = 32'hf9;
memory[3727] = 32'hfa;
memory[3728] = 32'hfb;
memory[3729] = 32'hfc;
memory[3730] = 32'hfd;
memory[3731] = 32'hfe;
memory[3732] = 32'he1;
memory[3733] = 32'he2;
memory[3734] = 32'he3;
memory[3735] = 32'he4;
memory[3736] = 32'he5;
memory[3737] = 32'he6;
memory[3738] = 32'he7;
memory[3739] = 32'he8;
memory[3740] = 32'he9;
memory[3741] = 32'hea;
memory[3742] = 32'heb;
memory[3743] = 32'hec;
memory[3744] = 32'hed;
memory[3745] = 32'hee;
memory[3746] = 32'hef;
memory[3747] = 32'hf0;
memory[3748] = 32'hf1;
memory[3749] = 32'hf2;
memory[3750] = 32'hf3;
memory[3751] = 32'hf4;
memory[3752] = 32'hf5;
memory[3753] = 32'hf6;
memory[3754] = 32'hf7;
memory[3755] = 32'hf8;
memory[3756] = 32'hf9;
memory[3757] = 32'hfa;
memory[3758] = 32'hfb;
memory[3759] = 32'hfc;
memory[3760] = 32'hfd;
memory[3761] = 32'hfe;
memory[3762] = 32'he1;
memory[3763] = 32'he2;
memory[3764] = 32'he3;
memory[3765] = 32'he4;
memory[3766] = 32'he5;
memory[3767] = 32'he6;
memory[3768] = 32'he7;
memory[3769] = 32'he8;
memory[3770] = 32'he9;
memory[3771] = 32'hea;
memory[3772] = 32'heb;
memory[3773] = 32'hec;
memory[3774] = 32'hed;
memory[3775] = 32'hf9;
memory[3776] = 32'hee;
memory[3777] = 32'heb;
memory[3778] = 32'hf0;
memory[3779] = 32'hfd;
memory[3780] = 32'hef;
memory[3781] = 32'he6;
memory[3782] = 32'he5;
memory[3783] = 32'hec;
memory[3784] = 32'hfb;
memory[3785] = 32'hfd;
memory[3786] = 32'hfe;
memory[3787] = 32'he1;
memory[3788] = 32'he2;
memory[3789] = 32'he3;
memory[3790] = 32'he4;
memory[3791] = 32'he5;
memory[3792] = 32'he6;
memory[3793] = 32'he7;
memory[3794] = 32'he8;
memory[3795] = 32'he9;
memory[3796] = 32'hea;
memory[3797] = 32'heb;
memory[3798] = 32'hec;
memory[3799] = 32'hed;
memory[3800] = 32'hee;
memory[3801] = 32'hef;
memory[3802] = 32'hf0;
memory[3803] = 32'hf1;
memory[3804] = 32'hf2;
memory[3805] = 32'hf3;
memory[3806] = 32'hf4;
memory[3807] = 32'hf5;
memory[3808] = 32'hf6;
memory[3809] = 32'hf7;
memory[3810] = 32'hf8;
memory[3811] = 32'hf9;
memory[3812] = 32'hfa;
memory[3813] = 32'hfb;
memory[3814] = 32'hfc;
memory[3815] = 32'hfd;
memory[3816] = 32'hfe;
memory[3817] = 32'he1;
memory[3818] = 32'he2;
memory[3819] = 32'he3;
memory[3820] = 32'he4;
memory[3821] = 32'he5;
memory[3822] = 32'he6;
memory[3823] = 32'he7;
memory[3824] = 32'he8;
memory[3825] = 32'he9;
memory[3826] = 32'hea;
memory[3827] = 32'heb;
memory[3828] = 32'hec;
memory[3829] = 32'hed;
memory[3830] = 32'hee;
memory[3831] = 32'hef;
memory[3832] = 32'hf0;
memory[3833] = 32'hf1;
memory[3834] = 32'hf2;
memory[3835] = 32'hf3;
memory[3836] = 32'hf4;
memory[3837] = 32'hf5;
memory[3838] = 32'hf6;
memory[3839] = 32'hf7;
memory[3840] = 32'hed;
memory[3841] = 32'hea;
memory[3842] = 32'hef;
memory[3843] = 32'hfc;
memory[3844] = 32'hf0;
memory[3845] = 32'he7;
memory[3846] = 32'he6;
memory[3847] = 32'hed;
memory[3848] = 32'hef;
memory[3849] = 32'hf0;
memory[3850] = 32'hf1;
memory[3851] = 32'hf2;
memory[3852] = 32'hf3;
memory[3853] = 32'hf4;
memory[3854] = 32'hf5;
memory[3855] = 32'hf6;
memory[3856] = 32'hf7;
memory[3857] = 32'hf8;
memory[3858] = 32'hf9;
memory[3859] = 32'hfa;
memory[3860] = 32'hfb;
memory[3861] = 32'hfc;
memory[3862] = 32'hfd;
memory[3863] = 32'hfe;
memory[3864] = 32'he1;
memory[3865] = 32'he2;
memory[3866] = 32'he3;
memory[3867] = 32'he4;
memory[3868] = 32'he5;
memory[3869] = 32'he6;
memory[3870] = 32'he7;
memory[3871] = 32'he8;
memory[3872] = 32'he9;
memory[3873] = 32'hea;
memory[3874] = 32'heb;
memory[3875] = 32'hec;
memory[3876] = 32'hed;
memory[3877] = 32'hee;
memory[3878] = 32'hef;
memory[3879] = 32'hf0;
memory[3880] = 32'hf1;
memory[3881] = 32'hf2;
memory[3882] = 32'hf3;
memory[3883] = 32'hf4;
memory[3884] = 32'hf5;
memory[3885] = 32'hf6;
memory[3886] = 32'hf7;
memory[3887] = 32'hf8;
memory[3888] = 32'hf9;
memory[3889] = 32'hfa;
memory[3890] = 32'hfb;
memory[3891] = 32'hfc;
memory[3892] = 32'hfd;
memory[3893] = 32'hfe;
memory[3894] = 32'he1;
memory[3895] = 32'he2;
memory[3896] = 32'he3;
memory[3897] = 32'he4;
memory[3898] = 32'he5;
memory[3899] = 32'he6;
memory[3900] = 32'he7;
memory[3901] = 32'he8;
memory[3902] = 32'he9;
memory[3903] = 32'hea;
memory[3904] = 32'heb;
memory[3905] = 32'he9;
memory[3906] = 32'hee;
memory[3907] = 32'hfb;
memory[3908] = 32'hf1;
memory[3909] = 32'he8;
memory[3910] = 32'he7;
memory[3911] = 32'he9;
memory[3912] = 32'hea;
memory[3913] = 32'heb;
memory[3914] = 32'hec;
memory[3915] = 32'hed;
memory[3916] = 32'hee;
memory[3917] = 32'hef;
memory[3918] = 32'hf0;
memory[3919] = 32'hf1;
memory[3920] = 32'hf2;
memory[3921] = 32'hf3;
memory[3922] = 32'hf4;
memory[3923] = 32'hf5;
memory[3924] = 32'hf6;
memory[3925] = 32'hf7;
memory[3926] = 32'hf8;
memory[3927] = 32'hf9;
memory[3928] = 32'hfa;
memory[3929] = 32'hfb;
memory[3930] = 32'hfc;
memory[3931] = 32'hfd;
memory[3932] = 32'hfe;
memory[3933] = 32'he1;
memory[3934] = 32'he2;
memory[3935] = 32'he3;
memory[3936] = 32'he4;
memory[3937] = 32'he5;
memory[3938] = 32'he6;
memory[3939] = 32'he7;
memory[3940] = 32'he8;
memory[3941] = 32'he9;
memory[3942] = 32'hea;
memory[3943] = 32'heb;
memory[3944] = 32'hec;
memory[3945] = 32'hed;
memory[3946] = 32'hee;
memory[3947] = 32'hef;
memory[3948] = 32'hf0;
memory[3949] = 32'hf1;
memory[3950] = 32'hf2;
memory[3951] = 32'hf3;
memory[3952] = 32'hf4;
memory[3953] = 32'hf5;
memory[3954] = 32'hf6;
memory[3955] = 32'hf7;
memory[3956] = 32'hf8;
memory[3957] = 32'hf9;
memory[3958] = 32'hfa;
memory[3959] = 32'hfb;
memory[3960] = 32'hfc;
memory[3961] = 32'hfd;
memory[3962] = 32'hfe;
memory[3963] = 32'he1;
memory[3964] = 32'he2;
memory[3965] = 32'he3;
memory[3966] = 32'he4;
memory[3967] = 32'he5;
memory[3968] = 32'he6;
memory[3969] = 32'he7;
memory[3970] = 32'hed;
memory[3971] = 32'hfa;
memory[3972] = 32'hf2;
memory[3973] = 32'he9;
memory[3974] = 32'heb;
memory[3975] = 32'hec;
memory[3976] = 32'hed;
memory[3977] = 32'hee;
memory[3978] = 32'hef;
memory[3979] = 32'hf0;
memory[3980] = 32'hf1;
memory[3981] = 32'hf2;
memory[3982] = 32'hf3;
memory[3983] = 32'hf4;
memory[3984] = 32'hf5;
memory[3985] = 32'hf6;
memory[3986] = 32'hf7;
memory[3987] = 32'hf8;
memory[3988] = 32'hf9;
memory[3989] = 32'hfa;
memory[3990] = 32'hfb;
memory[3991] = 32'hfc;
memory[3992] = 32'hfd;
memory[3993] = 32'hfe;
memory[3994] = 32'he1;
memory[3995] = 32'he2;
memory[3996] = 32'he3;
memory[3997] = 32'he4;
memory[3998] = 32'he5;
memory[3999] = 32'he6;
memory[4000] = 32'he7;
memory[4001] = 32'he8;
memory[4002] = 32'he9;
memory[4003] = 32'hea;
memory[4004] = 32'heb;
memory[4005] = 32'hec;
memory[4006] = 32'hed;
memory[4007] = 32'hee;
memory[4008] = 32'hef;
memory[4009] = 32'hf0;
memory[4010] = 32'hf1;
memory[4011] = 32'hf2;
memory[4012] = 32'hf3;
memory[4013] = 32'hf4;
memory[4014] = 32'hf5;
memory[4015] = 32'hf6;
memory[4016] = 32'hf7;
memory[4017] = 32'hf8;
memory[4018] = 32'hf9;
memory[4019] = 32'hfa;
memory[4020] = 32'hfb;
memory[4021] = 32'hfc;
memory[4022] = 32'hfd;
memory[4023] = 32'hfe;
memory[4024] = 32'he1;
memory[4025] = 32'he2;
memory[4026] = 32'he3;
memory[4027] = 32'he4;
memory[4028] = 32'he5;
memory[4029] = 32'he6;
memory[4030] = 32'he7;
memory[4031] = 32'he8;
memory[4032] = 32'he9;
memory[4033] = 32'hea;
memory[4034] = 32'heb;
memory[4035] = 32'hf9;
memory[4036] = 32'hf3;
memory[4037] = 32'hf5;
memory[4038] = 32'hf6;
memory[4039] = 32'hf7;
memory[4040] = 32'hf8;
memory[4041] = 32'hf9;
memory[4042] = 32'hfa;
memory[4043] = 32'hfb;
memory[4044] = 32'hfc;
memory[4045] = 32'hfd;
memory[4046] = 32'hfe;
memory[4047] = 32'he1;
memory[4048] = 32'he2;
memory[4049] = 32'he3;
memory[4050] = 32'he4;
memory[4051] = 32'he5;
memory[4052] = 32'he6;
memory[4053] = 32'he7;
memory[4054] = 32'he8;
memory[4055] = 32'he9;
memory[4056] = 32'hea;
memory[4057] = 32'heb;
memory[4058] = 32'hec;
memory[4059] = 32'hed;
memory[4060] = 32'hee;
memory[4061] = 32'hef;
memory[4062] = 32'hf0;
memory[4063] = 32'hf1;
memory[4064] = 32'hf2;
memory[4065] = 32'hf3;
memory[4066] = 32'hf4;
memory[4067] = 32'hf5;
memory[4068] = 32'hf6;
memory[4069] = 32'hf7;
memory[4070] = 32'hf8;
memory[4071] = 32'hf9;
memory[4072] = 32'hfa;
memory[4073] = 32'hfb;
memory[4074] = 32'hfc;
memory[4075] = 32'hfd;
memory[4076] = 32'hfe;
memory[4077] = 32'he1;
memory[4078] = 32'he2;
memory[4079] = 32'he3;
memory[4080] = 32'he4;
memory[4081] = 32'he5;
memory[4082] = 32'he6;
memory[4083] = 32'he7;
memory[4084] = 32'he8;
memory[4085] = 32'he9;
memory[4086] = 32'hea;
memory[4087] = 32'heb;
memory[4088] = 32'hec;
memory[4089] = 32'hed;
memory[4090] = 32'hee;
memory[4091] = 32'hef;
memory[4092] = 32'hf0;
memory[4093] = 32'hf1;
memory[4094] = 32'hf2;
memory[4095] = 32'hf3;
memory[4096] = 32'hf4;
memory[4097] = 32'hf5;
memory[4098] = 32'hf6;
memory[4099] = 32'hf7;
memory[4100] = 32'h63;
memory[4101] = 32'h63;
memory[4102] = 32'h63;
memory[4103] = 32'h63;
memory[4104] = 32'h63;
memory[4105] = 32'h63;
memory[4106] = 32'h63;
memory[4107] = 32'h63;
memory[4108] = 32'h63;
memory[4109] = 32'h63;
memory[4110] = 32'h63;
memory[4111] = 32'h63;
memory[4112] = 32'h63;
memory[4113] = 32'h63;
memory[4114] = 32'h63;
memory[4115] = 32'h63;
memory[4116] = 32'h0;




 
    end
   
    always @(posedge Clk) 
    begin
        if (MemWrite)   
        begin                           
//            if(whb == 2'b0)
//            begin
                memory[Address[15:2]] <= WriteData;
//            end
            
//            else if(whb == 2'b01)
//            begin
//                memory[Address[15:2]] <= {16'b0,WriteData[15:0]};
//            end
                
//            else if(whb == 2'b10)
//            begin
//                memory[Address[15:2]] <= {24'b0,WriteData[7:0]};
//            end
        end
    end
    
    always @(*) 
    begin
        if (MemRead)   
        begin                           
//            if(whb == 2'b0)
//            begin
                ReadData <= memory[Address[15:2]];
//            end
            
//            else if(whb == 2'b01)
//            begin
//                if(memory[Address[15:2]][15] == 0) begin
//                    ReadData <= {16'b0,memory[Address[15:2]][15:0]};
//                end
//                else begin
//                    ReadData <= {16'b1111111111111111,memory[Address[15:2]][15:0]};
//                end
//            end
                
//            else if(whb == 2'b10)
//            begin
//                if(memory[Address[11:2]][7] == 0) begin
//                    ReadData <= {24'b0,memory[Address[15:2]][7:0]};
//                end
//                else begin
//                    ReadData <= {24'b111111111111111111111111,memory[Address[15:2]][7:0]};
//                end
//            end
        end
    end
endmodule
